* Extracted by KLayout with SKY130 LVS runset on : 15/11/2024 23:50

.SUBCKT cap_vpp_04p4x04p6_l1m1m2_noshield SUB C1 C0
C$1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield
.ENDS cap_vpp_04p4x04p6_l1m1m2_noshield
