** sch_path: /Users/martin/Source/PEX-mjk/designs/nmos_diode/nmos_diode.sch
**.subckt nmos_diode VDD VSS
*.iopin VDD
*.iopin VSS
XM2 VDD VDD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
**** begin user architecture code


* .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt
* .op


**** end user architecture code
**.ends
.end
