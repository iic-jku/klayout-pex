* Extracted by KLayout with SKY130 LVS runset on : 08/11/2024 23:00

.SUBCKT sideoverlap_complex_li1_m1
.ENDS sideoverlap_complex_li1_m1
