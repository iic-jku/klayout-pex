* Extracted by KLayout with SKY130 LVS runset on : 07/11/2024 20:20

.SUBCKT sideoverlap_simple_plates_li1_m1
.ENDS sideoverlap_simple_plates_li1_m1
