* Extracted by KLayout with SKY130 LVS runset on : 18/10/2024 22:27

.SUBCKT sideoverlap_fingered_li1_m1
.ENDS sideoverlap_fingered_li1_m1
