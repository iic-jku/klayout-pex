sky130hs_lib.cdl