nmos_diode2.spice