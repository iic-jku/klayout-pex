* Extracted by KLayout with SKY130 LVS runset on : 08/11/2024 17:27

.SUBCKT sideoverlap_shielding_simple_plates_li1_m1_m2
.ENDS sideoverlap_shielding_simple_plates_li1_m1_m2
