* Extracted by KLayout with SKY130 LVS runset on : 09/10/2024 18:22

.SUBCKT single_plate_100um_x_100um_li1_over_substrate
.ENDS single_plate_100um_x_100um_li1_over_substrate
