* Extracted by KLayout with SKY130 LVS runset on : 13/09/2024 20:33

.SUBCKT cap_mim_m3_w18p9_l5p1
C$1 mimcap_bot mimcap_top sky130_fd_pr__model__cap_mim C=1.9278e-13 A=96.39 P=48
.ENDS cap_mim_m3_w18p9_l5p1
