nmos_diode.spice