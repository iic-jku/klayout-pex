* Extracted by KLayout on : 07/10/2024 17:06

.SUBCKT Contact
.ENDS Contact

.SUBCKT ntap
.ENDS ntap
