* Extracted by KLayout with SKY130 LVS runset on : 20/11/2024 15:49

.SUBCKT near_body_shield_li1_m1
.ENDS near_body_shield_li1_m1
