* Extracted by KLayout with SKY130 LVS runset on : 21/08/2024 18:01

.SUBCKT cap_vpp_04p4x04p6_l1m1m2_noshield
X1 C0 C1 SUB sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield
.ENDS cap_vpp_04p4x04p6_l1m1m2_noshield
