* Extracted by KLayout with SKY130 LVS runset on : 26/07/2024 16:19

.SUBCKT nmos_diode2
M$1 VDD VDD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 AS=0.126 AD=0.126
+ PS=1.44 PD=1.44
.ENDS nmos_diode2
