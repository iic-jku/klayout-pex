* Extracted by KLayout with SKY130 LVS runset on : 18/09/2024 19:04

.SUBCKT cap_mim_m3_w18p9_l5p1
C$1 \$1 \$2 sky130_fd_pr__model__cap_mim C=2.080738e-13 A=104.0369 P=49.23
.ENDS cap_mim_m3_w18p9_l5p1
