** sch_path: /Users/martin/Source/PEX-mjk/designs/nmos_diode2/nmos_diode2.sch
**.subckt nmos_diode2 VDD VSS
*.iopin VDD
*.iopin VSS
XM1 VDD VDD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 m=1
**** begin user architecture code


* .lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt
* .op


**** end user architecture code
**.ends
.end
