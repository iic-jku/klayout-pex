* Extracted by KLayout with SKY130 LVS runset on : 21/11/2024 17:38

.SUBCKT sidewall_net_uturn_l1_redux
.ENDS sidewall_net_uturn_l1_redux
