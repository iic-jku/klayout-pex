* Extracted by KLayout with SKY130 LVS runset on : 11/10/2024 17:32

.SUBCKT sidewall_100um_x_100um_distance_200nm_li1
.ENDS sidewall_100um_x_100um_distance_200nm_li1
