* Extracted by KLayout with SKY130 LVS runset on : 30/09/2024 15:36

.SUBCKT single_wire_met1_16x2
.ENDS single_wire_met1_16x2
