* Extracted by KLayout with SKY130 LVS runset on : 24/10/2024 22:11

.SUBCKT sideoverlap_plates_li1_m1
.ENDS sideoverlap_plates_li1_m1
