* Extracted by KLayout with SKY130 LVS runset on : 21/06/2024 21:30

.SUBCKT nmos_diode
M$1 VDD VDD VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 AS=0.84 AD=0.84 PS=6.56
+ PD=6.56
.ENDS nmos_diode
