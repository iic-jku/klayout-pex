* Extracted by KLayout on : 09/10/2024 17:13

.SUBCKT sky130_fd_sc_hs__a2111o_1 VGND B1 C1 A1 X A2 D1 VPWR VPB VNB
M$1 X \$7 VPWR VPB pfet_01v8 L=150000U W=1120000U AS=308000000000P
+ AD=308000000000P PS=2790000U PD=2790000U
M$2 VPWR A1 \$11 VPB pfet_01v8 L=150000U W=1000000U AS=275000000000P
+ AD=170000000000P PS=2550000U PD=1340000U
M$3 \$11 A2 VPWR VPB pfet_01v8 L=150000U W=1000000U AS=170000000000P
+ AD=150000000000P PS=1340000U PD=1300000U
M$4 \$14 B1 \$11 VPB pfet_01v8 L=150000U W=1000000U AS=150000000000P
+ AD=120000000000P PS=1300000U PD=1240000U
M$5 \$15 C1 \$14 VPB pfet_01v8 L=150000U W=1000000U AS=120000000000P
+ AD=120000000000P PS=1240000U PD=1240000U
M$6 \$7 D1 \$15 VPB pfet_01v8 L=150000U W=1000000U AS=120000000000P
+ AD=275000000000P PS=1240000U PD=2550000U
M$7 \$8 A1 \$7 VNB nfet_01v8_lvt L=150000U W=640000U AS=169600000000P
+ AD=67200000000P PS=1810000U PD=850000U
M$8 VGND A2 \$8 VNB nfet_01v8_lvt L=150000U W=640000U AS=67200000000P
+ AD=124800000000P PS=850000U PD=1030000U
M$9 \$7 B1 VGND VNB nfet_01v8_lvt L=150000U W=640000U AS=124800000000P
+ AD=89600000000P PS=1030000U PD=920000U
M$10 VGND C1 \$7 VNB nfet_01v8_lvt L=150000U W=640000U AS=89600000000P
+ AD=150400000000P PS=920000U PD=1110000U
M$11 \$7 D1 VGND VNB nfet_01v8_lvt L=150000U W=640000U AS=150400000000P
+ AD=169600000000P PS=1110000U PD=1810000U
M$12 X \$7 VGND VNB nfet_01v8_lvt L=150000U W=740000U AS=196100000000P
+ AD=196100000000P PS=2010000U PD=2010000U
CCext31 0 \$11 8.10039e-17 PEX_CAP
CCext41 A1 \$11 3.91575e-16 PEX_CAP
CCext51 A2 \$11 2.2824e-16 PEX_CAP
CCext61 B1 \$11 3.33861e-16 PEX_CAP
CCext101 VPWR \$11 2.01302e-16 PEX_CAP
CCext11 \$11 0 5.26785162e-16 PEX_CAP
CCext32 0 \$7 2.65253e-16 PEX_CAP
CCext42 A1 \$7 2.23253e-16 PEX_CAP
CCext52 A2 \$7 9.53683e-17 PEX_CAP
CCext62 B1 \$7 1.7429e-16 PEX_CAP
CCext72 C1 \$7 1.04e-16 PEX_CAP
CCext82 D1 \$7 4.01133e-16 PEX_CAP
CCext92 VGND \$7 3.71912e-16 PEX_CAP
CCext102 VPWR \$7 3.75257e-16 PEX_CAP
CCext112 X \$7 4.06551e-16 PEX_CAP
CCext22 \$7 0 1.7328961e-15 PEX_CAP
CCext43 A1 0 2.86244e-16 PEX_CAP
CCext53 A2 0 8.79653e-17 PEX_CAP
CCext63 B1 0 2.19135e-16 PEX_CAP
CCext73 C1 0 1.25201e-16 PEX_CAP
CCext83 D1 0 1.18603e-16 PEX_CAP
CCext93 VGND 0 1.35941e-16 PEX_CAP
CCext103 VPWR 0 1.51499e-16 PEX_CAP
CCext113 X 0 8.59454e-17 PEX_CAP
CCext54 A2 A1 1.18505e-16 PEX_CAP
CCext94 VGND A1 1.08337e-16 PEX_CAP
CCext104 VPWR A1 1.2477e-16 PEX_CAP
CCext44 A1 0 3.62983917e-16 PEX_CAP
CCext65 B1 A2 1.32528e-16 PEX_CAP
CCext95 VGND A2 9.22956e-17 PEX_CAP
CCext105 VPWR A2 1.30159e-16 PEX_CAP
CCext76 C1 B1 1.6494e-16 PEX_CAP
CCext96 VGND B1 1.42284e-16 PEX_CAP
CCext66 B1 0 3.37011557e-16 PEX_CAP
CCext87 D1 C1 1.10351e-16 PEX_CAP
CCext97 VGND C1 1.28679e-16 PEX_CAP
CCext98 VGND D1 9.34773e-17 PEX_CAP
CCext119 X VGND 1.05534e-16 PEX_CAP
CCext1110 X VPWR 1.27279e-16 PEX_CAP
.ENDS sky130_fd_sc_hs__a2111o_1
