* Extracted by KLayout with SKY130 LVS runset on : 11/10/2024 20:41

.SUBCKT overlap_plates_100um_x_100um_li1_m1
.ENDS overlap_plates_100um_x_100um_li1_m1
