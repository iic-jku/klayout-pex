.subckt cap_mim_m3_w18p9_l5p1
C1 mimcap_bot mimcap_top sky130_fd_pr__model__cap_mim C=1.9278e-13 A=96.39 P=48
.ends cap_mim_m3_w18p9_l5p1
