* Extracted by KLayout with SKY130 LVS runset on : 15/10/2024 20:44

.SUBCKT overlap_plates_100um_x_100um_li1_m1_m2_m3
.ENDS overlap_plates_100um_x_100um_li1_m1_m2_m3
