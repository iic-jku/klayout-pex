* Extracted by KLayout with SKY130 LVS runset on : 21/11/2024 16:25

.SUBCKT sidewall_cap_vpp_04p4x04p6_l1_redux
.ENDS sidewall_cap_vpp_04p4x04p6_l1_redux
