* Extracted by KLayout with SKY130 LVS runset on : 22/10/2024 16:25

.SUBCKT sideoverlap_fingered_li1_m1_patternA
.ENDS sideoverlap_fingered_li1_m1_patternA
