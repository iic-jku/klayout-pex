.subckt single_wire_met1_16x2
.ends single_wire_met1_16x2
