* NGSPICE file created from gcd.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt gcd VGND VPWR clk operands_bits_A[0] operands_bits_A[100] operands_bits_A[101]
+ operands_bits_A[102] operands_bits_A[103] operands_bits_A[104] operands_bits_A[105]
+ operands_bits_A[106] operands_bits_A[107] operands_bits_A[108] operands_bits_A[109]
+ operands_bits_A[10] operands_bits_A[110] operands_bits_A[111] operands_bits_A[112]
+ operands_bits_A[113] operands_bits_A[114] operands_bits_A[115] operands_bits_A[116]
+ operands_bits_A[117] operands_bits_A[118] operands_bits_A[119] operands_bits_A[11]
+ operands_bits_A[120] operands_bits_A[121] operands_bits_A[122] operands_bits_A[123]
+ operands_bits_A[124] operands_bits_A[125] operands_bits_A[126] operands_bits_A[127]
+ operands_bits_A[12] operands_bits_A[13] operands_bits_A[14] operands_bits_A[15]
+ operands_bits_A[16] operands_bits_A[17] operands_bits_A[18] operands_bits_A[19]
+ operands_bits_A[1] operands_bits_A[20] operands_bits_A[21] operands_bits_A[22] operands_bits_A[23]
+ operands_bits_A[24] operands_bits_A[25] operands_bits_A[26] operands_bits_A[27]
+ operands_bits_A[28] operands_bits_A[29] operands_bits_A[2] operands_bits_A[30] operands_bits_A[31]
+ operands_bits_A[32] operands_bits_A[33] operands_bits_A[34] operands_bits_A[35]
+ operands_bits_A[36] operands_bits_A[37] operands_bits_A[38] operands_bits_A[39]
+ operands_bits_A[3] operands_bits_A[40] operands_bits_A[41] operands_bits_A[42] operands_bits_A[43]
+ operands_bits_A[44] operands_bits_A[45] operands_bits_A[46] operands_bits_A[47]
+ operands_bits_A[48] operands_bits_A[49] operands_bits_A[4] operands_bits_A[50] operands_bits_A[51]
+ operands_bits_A[52] operands_bits_A[53] operands_bits_A[54] operands_bits_A[55]
+ operands_bits_A[56] operands_bits_A[57] operands_bits_A[58] operands_bits_A[59]
+ operands_bits_A[5] operands_bits_A[60] operands_bits_A[61] operands_bits_A[62] operands_bits_A[63]
+ operands_bits_A[64] operands_bits_A[65] operands_bits_A[66] operands_bits_A[67]
+ operands_bits_A[68] operands_bits_A[69] operands_bits_A[6] operands_bits_A[70] operands_bits_A[71]
+ operands_bits_A[72] operands_bits_A[73] operands_bits_A[74] operands_bits_A[75]
+ operands_bits_A[76] operands_bits_A[77] operands_bits_A[78] operands_bits_A[79]
+ operands_bits_A[7] operands_bits_A[80] operands_bits_A[81] operands_bits_A[82] operands_bits_A[83]
+ operands_bits_A[84] operands_bits_A[85] operands_bits_A[86] operands_bits_A[87]
+ operands_bits_A[88] operands_bits_A[89] operands_bits_A[8] operands_bits_A[90] operands_bits_A[91]
+ operands_bits_A[92] operands_bits_A[93] operands_bits_A[94] operands_bits_A[95]
+ operands_bits_A[96] operands_bits_A[97] operands_bits_A[98] operands_bits_A[99]
+ operands_bits_A[9] operands_bits_B[0] operands_bits_B[100] operands_bits_B[101]
+ operands_bits_B[102] operands_bits_B[103] operands_bits_B[104] operands_bits_B[105]
+ operands_bits_B[106] operands_bits_B[107] operands_bits_B[108] operands_bits_B[109]
+ operands_bits_B[10] operands_bits_B[110] operands_bits_B[111] operands_bits_B[112]
+ operands_bits_B[113] operands_bits_B[114] operands_bits_B[115] operands_bits_B[116]
+ operands_bits_B[117] operands_bits_B[118] operands_bits_B[119] operands_bits_B[11]
+ operands_bits_B[120] operands_bits_B[121] operands_bits_B[122] operands_bits_B[123]
+ operands_bits_B[124] operands_bits_B[125] operands_bits_B[126] operands_bits_B[127]
+ operands_bits_B[12] operands_bits_B[13] operands_bits_B[14] operands_bits_B[15]
+ operands_bits_B[16] operands_bits_B[17] operands_bits_B[18] operands_bits_B[19]
+ operands_bits_B[1] operands_bits_B[20] operands_bits_B[21] operands_bits_B[22] operands_bits_B[23]
+ operands_bits_B[24] operands_bits_B[25] operands_bits_B[26] operands_bits_B[27]
+ operands_bits_B[28] operands_bits_B[29] operands_bits_B[2] operands_bits_B[30] operands_bits_B[31]
+ operands_bits_B[32] operands_bits_B[33] operands_bits_B[34] operands_bits_B[35]
+ operands_bits_B[36] operands_bits_B[37] operands_bits_B[38] operands_bits_B[39]
+ operands_bits_B[3] operands_bits_B[40] operands_bits_B[41] operands_bits_B[42] operands_bits_B[43]
+ operands_bits_B[44] operands_bits_B[45] operands_bits_B[46] operands_bits_B[47]
+ operands_bits_B[48] operands_bits_B[49] operands_bits_B[4] operands_bits_B[50] operands_bits_B[51]
+ operands_bits_B[52] operands_bits_B[53] operands_bits_B[54] operands_bits_B[55]
+ operands_bits_B[56] operands_bits_B[57] operands_bits_B[58] operands_bits_B[59]
+ operands_bits_B[5] operands_bits_B[60] operands_bits_B[61] operands_bits_B[62] operands_bits_B[63]
+ operands_bits_B[64] operands_bits_B[65] operands_bits_B[66] operands_bits_B[67]
+ operands_bits_B[68] operands_bits_B[69] operands_bits_B[6] operands_bits_B[70] operands_bits_B[71]
+ operands_bits_B[72] operands_bits_B[73] operands_bits_B[74] operands_bits_B[75]
+ operands_bits_B[76] operands_bits_B[77] operands_bits_B[78] operands_bits_B[79]
+ operands_bits_B[7] operands_bits_B[80] operands_bits_B[81] operands_bits_B[82] operands_bits_B[83]
+ operands_bits_B[84] operands_bits_B[85] operands_bits_B[86] operands_bits_B[87]
+ operands_bits_B[88] operands_bits_B[89] operands_bits_B[8] operands_bits_B[90] operands_bits_B[91]
+ operands_bits_B[92] operands_bits_B[93] operands_bits_B[94] operands_bits_B[95]
+ operands_bits_B[96] operands_bits_B[97] operands_bits_B[98] operands_bits_B[99]
+ operands_bits_B[9] operands_rdy operands_val reset result_bits_data[0] result_bits_data[100]
+ result_bits_data[101] result_bits_data[102] result_bits_data[103] result_bits_data[104]
+ result_bits_data[105] result_bits_data[106] result_bits_data[107] result_bits_data[108]
+ result_bits_data[109] result_bits_data[10] result_bits_data[110] result_bits_data[111]
+ result_bits_data[112] result_bits_data[113] result_bits_data[114] result_bits_data[115]
+ result_bits_data[116] result_bits_data[117] result_bits_data[118] result_bits_data[119]
+ result_bits_data[11] result_bits_data[120] result_bits_data[121] result_bits_data[122]
+ result_bits_data[123] result_bits_data[124] result_bits_data[125] result_bits_data[126]
+ result_bits_data[127] result_bits_data[12] result_bits_data[13] result_bits_data[14]
+ result_bits_data[15] result_bits_data[16] result_bits_data[17] result_bits_data[18]
+ result_bits_data[19] result_bits_data[1] result_bits_data[20] result_bits_data[21]
+ result_bits_data[22] result_bits_data[23] result_bits_data[24] result_bits_data[25]
+ result_bits_data[26] result_bits_data[27] result_bits_data[28] result_bits_data[29]
+ result_bits_data[2] result_bits_data[30] result_bits_data[31] result_bits_data[32]
+ result_bits_data[33] result_bits_data[34] result_bits_data[35] result_bits_data[36]
+ result_bits_data[37] result_bits_data[38] result_bits_data[39] result_bits_data[3]
+ result_bits_data[40] result_bits_data[41] result_bits_data[42] result_bits_data[43]
+ result_bits_data[44] result_bits_data[45] result_bits_data[46] result_bits_data[47]
+ result_bits_data[48] result_bits_data[49] result_bits_data[4] result_bits_data[50]
+ result_bits_data[51] result_bits_data[52] result_bits_data[53] result_bits_data[54]
+ result_bits_data[55] result_bits_data[56] result_bits_data[57] result_bits_data[58]
+ result_bits_data[59] result_bits_data[5] result_bits_data[60] result_bits_data[61]
+ result_bits_data[62] result_bits_data[63] result_bits_data[64] result_bits_data[65]
+ result_bits_data[66] result_bits_data[67] result_bits_data[68] result_bits_data[69]
+ result_bits_data[6] result_bits_data[70] result_bits_data[71] result_bits_data[72]
+ result_bits_data[73] result_bits_data[74] result_bits_data[75] result_bits_data[76]
+ result_bits_data[77] result_bits_data[78] result_bits_data[79] result_bits_data[7]
+ result_bits_data[80] result_bits_data[81] result_bits_data[82] result_bits_data[83]
+ result_bits_data[84] result_bits_data[85] result_bits_data[86] result_bits_data[87]
+ result_bits_data[88] result_bits_data[89] result_bits_data[8] result_bits_data[90]
+ result_bits_data[91] result_bits_data[92] result_bits_data[93] result_bits_data[94]
+ result_bits_data[95] result_bits_data[96] result_bits_data[97] result_bits_data[98]
+ result_bits_data[99] result_bits_data[9] result_rdy result_val
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3155_ _1194_ _1203_ _1205_ _0779_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3086_ net283 GCDdpath0.B_reg\[120\] VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3988_ _0643_ _0701_ _1938_ _0644_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__o31a_1
XFILLER_0_162_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2939_ _0913_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4609_ _2405_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4960_ clknet_leaf_34_clk _0292_ _0036_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3911_ net61 _1804_ _1734_ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__or3_1
X_4891_ _2457_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3842_ _1770_ _0837_ _1722_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3773_ _1748_ _1754_ _1326_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_172_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2724_ _0773_ _0774_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2655_ _0660_ _0700_ _0662_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_112_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2586_ net293 _0636_ GCDdpath0.B_reg\[15\] _0635_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_160_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4325_ _2206_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_35_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4256_ _2082_ VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__buf_2
X_3207_ _1158_ _1257_ _1149_ _1140_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__or4_1
X_4187_ GCDdpath0.B_reg\[126\] net158 _1904_ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__mux2_1
X_3138_ net392 _0840_ _0842_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3069_ _1111_ _1113_ _1112_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_164_Left_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_Left_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4110_ _0620_ _0630_ _2016_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__nand3_1
X_5090_ clknet_leaf_32_clk _0422_ _0166_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4041_ net41 _1983_ _1984_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4943_ clknet_leaf_43_clk _0275_ _0019_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4874_ _2455_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3825_ net334 _1793_ _1798_ _1559_ _1799_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__o221a_1
XFILLER_0_144_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3756_ _1740_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2707_ _0738_ _0744_ _0751_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__nor4_1
XFILLER_0_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3687_ net97 _1583_ _1517_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__o21a_1
X_2638_ _0686_ _0687_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput264 net264 VGND VGND VPWR VPWR result_bits_data[103] sky130_fd_sc_hd__clkbuf_4
X_2569_ net282 GCDdpath0.B_reg\[11\] VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__xor2_1
Xoutput275 net275 VGND VGND VPWR VPWR result_bits_data[113] sky130_fd_sc_hd__clkbuf_4
Xoutput286 net286 VGND VGND VPWR VPWR result_bits_data[123] sky130_fd_sc_hd__clkbuf_4
Xoutput297 net297 VGND VGND VPWR VPWR result_bits_data[18] sky130_fd_sc_hd__clkbuf_4
X_4308_ _2194_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4239_ GCDdpath0.B_reg\[111\] net142 _2142_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3610_ _1405_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4590_ net365 _2392_ _2386_ VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3541_ net119 _1432_ _1479_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3472_ _1405_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5142_ clknet_leaf_12_clk _0474_ _0218_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dfrtp_4
X_5073_ clknet_leaf_44_clk _0405_ _0149_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dfrtp_4
X_4024_ net303 _1970_ _1911_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4926_ clknet_leaf_39_clk _0002_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_158_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4857_ _2451_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3808_ _1784_ _1774_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4788_ _2441_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3739_ _0725_ _1725_ _1187_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2972_ GCDdpath0.B_reg\[105\] net266 VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _2428_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4642_ _2416_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4573_ net291 _2380_ _2372_ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3524_ _0861_ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3455_ _1060_ _1475_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3386_ _0977_ _0999_ _1016_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__nand3_2
X_5125_ clknet_leaf_21_clk _0457_ _0201_ VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5056_ clknet_leaf_40_clk _0388_ _0132_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4007_ _0655_ _1915_ VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4909_ _2460_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _0570_ _0515_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3171_ net358 GCDdpath0.B_reg\[73\] VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__or2b_1
XFILLER_0_174_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ _1005_ _0903_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2886_ _0935_ _0936_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4625_ _2414_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4556_ net296 _2368_ _2358_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3507_ _0808_ _0848_ _0976_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__a21o_1
X_4487_ net319 _2320_ _2316_ VGND VGND VPWR VPWR _2321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3438_ GCDdpath0.B_reg\[104\] _1464_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _1404_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__clkbuf_2
X_5108_ clknet_leaf_14_clk _0440_ _0184_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5039_ clknet_leaf_3_clk _0371_ _0115_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput120 operands_bits_A[92] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
Xinput131 operands_bits_B[101] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_1
Xinput142 operands_bits_B[111] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xinput153 operands_bits_B[121] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xinput164 operands_bits_B[16] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_1
Xinput175 operands_bits_B[26] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_2
Xinput186 operands_bits_B[36] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_1
XFILLER_0_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput197 operands_bits_B[46] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ _0789_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2671_ _0720_ _0721_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4410_ GCDdpath0.B_reg\[60\] net213 _2256_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4341_ net367 _2217_ _2215_ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4272_ net262 _2168_ _2158_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3223_ _1156_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3154_ _1204_ GCDdpath0.B_reg\[42\] _0781_ _0780_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3085_ GCDdpath0.B_reg\[121\] net284 VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3987_ _0655_ _1915_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2938_ _0919_ _0920_ _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__or3b_1
XFILLER_0_115_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2869_ net358 GCDdpath0.B_reg\[73\] VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4608_ net299 _2404_ _2044_ VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4539_ GCDdpath0.B_reg\[22\] net171 _2356_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3910_ GCDdpath0.B_reg\[39\] _1872_ _1797_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4890_ _2457_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3841_ _1813_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3772_ _0710_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2723_ net326 GCDdpath0.B_reg\[44\] VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__or2b_1
XFILLER_0_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2654_ _0642_ _0702_ _0704_ _0639_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2585_ _0635_ GCDdpath0.B_reg\[15\] GCDdpath0.B_reg\[14\] VGND VGND VPWR VPWR _0636_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4324_ net372 _2205_ _2201_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4255_ GCDdpath0.B_reg\[106\] net136 _2156_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3206_ _1153_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__inv_2
X_4186_ _2108_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_1
X_3137_ _0712_ _0715_ _0716_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__o21bai_1
X_3068_ _1106_ _1108_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4040_ _1286_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4942_ clknet_leaf_45_clk _0274_ _0018_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4873_ _2454_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3824_ net75 _1506_ _1734_ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_31_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3755_ net345 _1739_ _1687_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2706_ _0752_ _0753_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__or3_1
XFILLER_0_160_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3686_ net395 _1296_ _1679_ _1680_ _1536_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ GCDdpath0.B_reg\[19\] net298 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ _0617_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__nand2_1
Xoutput265 net265 VGND VGND VPWR VPWR result_bits_data[104] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput276 net276 VGND VGND VPWR VPWR result_bits_data[114] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput287 net287 VGND VGND VPWR VPWR result_bits_data[124] sky130_fd_sc_hd__clkbuf_4
Xoutput298 net298 VGND VGND VPWR VPWR result_bits_data[19] sky130_fd_sc_hd__clkbuf_4
X_4307_ net378 _2193_ _2187_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__mux2_1
X_2499_ GCDdpath0.B_reg\[103\] GCDdpath0.B_reg\[102\] GCDdpath0.B_reg\[101\] GCDdpath0.B_reg\[100\]
+ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4238_ _2145_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _0584_ _0579_ _0582_ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3540_ GCDdpath0.B_reg\[91\] _1285_ _1549_ _1554_ _1536_ VGND VGND VPWR VPWR _1555_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3471_ _1494_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5141_ clknet_leaf_12_clk _0473_ _0217_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ clknet_leaf_44_clk _0404_ _0148_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4023_ net44 _1969_ _1898_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4925_ clknet_leaf_39_clk _0001_ VGND VGND VPWR VPWR GCDctrl0.state\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4856_ _2451_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3807_ _0752_ _0753_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4787_ _2440_ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3738_ _0718_ _1724_ _0844_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_144_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ net99 _1664_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_170_Right_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2971_ _1017_ _1018_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4710_ _2428_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641_ _2416_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4572_ GCDdpath0.B_reg\[12\] net160 _2370_ VGND VGND VPWR VPWR _2380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3523_ _0857_ _1529_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3454_ net264 _1445_ _1478_ _1480_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3385_ _1069_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__inv_2
X_5124_ clknet_leaf_14_clk _0456_ _0200_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dfrtp_4
X_5055_ clknet_leaf_1_clk _0387_ _0131_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_49_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
X_4006_ _1509_ _1950_ _1953_ _1954_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4908_ _2454_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4839_ _2449_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_6 net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _0914_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2954_ net366 _0895_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_106_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2885_ net363 GCDdpath0.B_reg\[78\] VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4624_ _2414_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4555_ GCDdpath0.B_reg\[17\] net165 _2356_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3506_ _0857_ _0860_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4486_ GCDdpath0.B_reg\[38\] net188 _2314_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3437_ _1027_ _1422_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_115_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ net257 net259 VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5107_ clknet_leaf_27_clk _0439_ _0183_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dfrtp_4
X_3299_ _1135_ _1136_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__nor2_1
X_5038_ clknet_leaf_7_clk _0370_ _0114_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput110 operands_bits_A[83] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xinput121 operands_bits_A[93] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xinput132 operands_bits_B[102] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput143 operands_bits_B[112] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
Xinput154 operands_bits_B[122] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xinput165 operands_bits_B[17] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
Xinput176 operands_bits_B[27] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput187 operands_bits_B[37] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
Xinput198 operands_bits_B[47] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2670_ net346 GCDdpath0.B_reg\[62\] VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4340_ GCDdpath0.B_reg\[81\] net236 _2213_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4271_ GCDdpath0.B_reg\[101\] net131 _2156_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3222_ _1270_ _1271_ _1272_ _0575_ _1157_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3153_ net324 VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3084_ net284 GCDdpath0.B_reg\[121\] VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3986_ _1937_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2937_ _0921_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2868_ _0915_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ GCDdpath0.B_reg\[1\] net168 _1495_ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2799_ GCDdpath0.B_reg\[95\] net382 VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4538_ _2313_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4469_ net398 _2307_ _2301_ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_171_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3840_ net331 _1812_ _1745_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3771_ _0839_ _1747_ _0715_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2722_ GCDdpath0.B_reg\[44\] net326 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2653_ _0640_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2584_ net294 VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4323_ GCDdpath0.B_reg\[86\] net241 _2199_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4254_ _2141_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3205_ _1070_ _1241_ _1249_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o211a_1
X_4185_ net290 _2107_ _1282_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__mux2_1
X_3136_ GCDdpath0.B_reg\[60\] net344 VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3067_ _1071_ _1092_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3969_ _1923_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_166_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4941_ clknet_leaf_45_clk _0273_ _0017_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4872_ reset VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3823_ GCDdpath0.B_reg\[51\] _1796_ _1797_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3754_ net86 _1738_ _1718_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2705_ _0754_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__or2_1
X_3685_ _0959_ _0964_ _1678_ _1326_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2636_ net298 GCDdpath0.B_reg\[19\] VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2567_ net292 GCDdpath0.B_reg\[13\] VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__xnor2_1
Xoutput266 net266 VGND VGND VPWR VPWR result_bits_data[105] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput277 net277 VGND VGND VPWR VPWR result_bits_data[115] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4306_ GCDdpath0.B_reg\[91\] net247 _2184_ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__mux2_1
Xoutput288 net288 VGND VGND VPWR VPWR result_bits_data[125] sky130_fd_sc_hd__clkbuf_4
Xoutput299 net299 VGND VGND VPWR VPWR result_bits_data[1] sky130_fd_sc_hd__clkbuf_4
X_2498_ _0544_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4237_ net274 _2143_ _2144_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__mux2_1
X_4168_ _2094_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3119_ _1169_ GCDdpath0.B_reg\[26\] _0639_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4099_ _2034_ _2035_ _1609_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3470_ net261 _1493_ _1489_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ clknet_leaf_13_clk _0472_ _0216_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dfrtp_4
X_5071_ clknet_leaf_43_clk _0403_ _0147_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dfrtp_4
X_4022_ GCDdpath0.B_reg\[23\] _1968_ _1892_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4924_ clknet_leaf_39_clk _0000_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_87_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4855_ _2451_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3806_ _1783_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_1
X_4786_ reset VGND VGND VPWR VPWR _2440_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_117_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3737_ net391 _1723_ _0816_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3668_ _1336_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2619_ GCDdpath0.B_reg\[21\] net301 VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3599_ _0901_ _1604_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2970_ _1019_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _2416_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4571_ _2379_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3522_ _1292_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3453_ net5 _1432_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3384_ _1029_ _1030_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__nor2_1
X_5123_ clknet_leaf_22_clk _0455_ _0199_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5054_ clknet_leaf_2_clk _0386_ _0130_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4005_ GCDdpath0.B_reg\[25\] _1516_ _1353_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4907_ _2459_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4838_ _2449_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4769_ _2437_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_168_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2953_ net367 GCDdpath0.B_reg\[81\] VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2884_ GCDdpath0.B_reg\[78\] net363 VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4623_ _2414_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4554_ _2367_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3505_ _1524_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4485_ _2319_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3436_ _1299_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _1403_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_1
X_5106_ clknet_leaf_30_clk _0438_ _0182_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3298_ _1299_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__buf_2
X_5037_ clknet_leaf_3_clk _0369_ _0113_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput100 operands_bits_A[74] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_1
Xinput111 operands_bits_A[84] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_1
Xinput122 operands_bits_A[94] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
Xinput133 operands_bits_B[103] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xinput144 operands_bits_B[113] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xinput155 operands_bits_B[123] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xinput166 operands_bits_B[18] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
Xinput177 operands_bits_B[28] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_1
XFILLER_0_99_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput188 operands_bits_B[38] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
XFILLER_0_37_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput199 operands_bits_B[48] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4270_ _2167_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_169_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3221_ _1152_ _1145_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3152_ _0794_ _1198_ _1201_ _1202_ _0792_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a41o_1
XFILLER_0_20_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3083_ _1130_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3985_ net308 _1936_ _1911_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2936_ GCDdpath0.B_reg\[72\] net357 VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2867_ _0916_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4606_ _2403_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2798_ net382 GCDdpath0.B_reg\[95\] VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__or2b_1
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4537_ _2355_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4468_ GCDdpath0.B_reg\[43\] net194 _2299_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__mux2_1
X_3419_ _1446_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4399_ net348 _2257_ _2258_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_165_Right_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3770_ net83 _1415_ _0517_ _1752_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__o31a_1
XFILLER_0_156_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2721_ _0770_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2652_ GCDdpath0.B_reg\[26\] net306 VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2583_ _0626_ _0627_ _0633_ _0619_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__o2bb2a_1
X_4322_ _2204_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4253_ _2155_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3204_ _1081_ _1254_ _1030_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__a21oi_1
X_4184_ GCDdpath0.B_reg\[127\] net159 _1904_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__mux2_1
X_3135_ GCDdpath0.B_reg\[61\] net345 VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3066_ _1098_ _1104_ _1110_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3968_ net312 _1922_ _1911_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2919_ net352 GCDdpath0.B_reg\[68\] VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__or2b_2
XFILLER_0_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3899_ _0791_ _1823_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_142_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ clknet_leaf_45_clk _0272_ _0016_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4871_ _2453_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3822_ _1295_ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3753_ GCDdpath0.B_reg\[61\] _1737_ _1684_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2704_ GCDdpath0.B_reg\[52\] net335 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3684_ _0959_ _1678_ _0964_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__a21oi_1
X_2635_ GCDdpath0.B_reg\[18\] net297 VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2566_ _0615_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput267 net267 VGND VGND VPWR VPWR result_bits_data[106] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4305_ _2192_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__clkbuf_1
Xoutput278 net278 VGND VGND VPWR VPWR result_bits_data[116] sky130_fd_sc_hd__clkbuf_4
Xoutput289 net289 VGND VGND VPWR VPWR result_bits_data[126] sky130_fd_sc_hd__clkbuf_4
X_2497_ _0545_ _0546_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_160_Left_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4236_ _2082_ VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4167_ net321 _2093_ _2041_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__mux2_1
X_3118_ net306 VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4098_ net292 net33 _1904_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__mux2_1
X_3049_ net279 GCDdpath0.B_reg\[117\] VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__and2b_1
XFILLER_0_167_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5070_ clknet_leaf_45_clk _0402_ _0146_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dfrtp_4
X_4021_ _0667_ _1967_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4923_ _2409_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4854_ _2451_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3805_ net337 _1782_ _1745_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4785_ _2439_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3736_ _0837_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3667_ GCDdpath0.B_reg\[73\] _1663_ _1598_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2618_ net301 GCDdpath0.B_reg\[21\] VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3598_ _0901_ _1604_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2549_ _0592_ _0595_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__and2b_1
X_4219_ net279 _2131_ _2129_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ net292 _2378_ _2372_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3521_ net381 _1445_ _1537_ _1538_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__o22a_1
XFILLER_0_170_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3452_ _0572_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3383_ _1326_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__buf_2
XFILLER_0_23_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5122_ clknet_leaf_22_clk _0454_ _0198_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5053_ clknet_leaf_39_clk _0385_ _0129_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4004_ _1951_ _1952_ _1511_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4906_ _2459_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4837_ _2447_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4768_ _2437_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3719_ net350 _1708_ _1687_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__mux2_1
X_4699_ _2425_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2952_ _0899_ _0907_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2883_ _0932_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4622_ _2413_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4553_ net297 _2366_ _2358_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3504_ net383 _1523_ _1489_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4484_ net320 _2318_ _2316_ VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3435_ _1463_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3366_ net275 _1402_ _1393_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5105_ clknet_leaf_30_clk _0437_ _0181_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dfrtp_4
X_3297_ _0517_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__clkbuf_2
X_5036_ clknet_leaf_3_clk _0368_ _0112_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput101 operands_bits_A[75] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xinput112 operands_bits_A[85] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
Xinput123 operands_bits_A[95] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xinput134 operands_bits_B[104] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
Xinput145 operands_bits_B[114] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_1
Xinput156 operands_bits_B[124] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_2
Xinput167 operands_bits_B[19] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_1
Xinput178 operands_bits_B[29] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_1
XFILLER_0_76_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput189 operands_bits_B[39] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__buf_1
XFILLER_0_99_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3220_ _0577_ _1146_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3151_ net319 _0793_ GCDdpath0.B_reg\[38\] VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3082_ _1131_ _1132_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3984_ net49 _1935_ _1898_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2935_ _0959_ _0962_ _0965_ _0984_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_28_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2866_ GCDdpath0.B_reg\[74\] net359 VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__or2b_1
XFILLER_0_115_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4605_ net310 _2402_ _2044_ VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2797_ _0731_ _0816_ _0846_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__o211a_2
XFILLER_0_142_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4536_ net303 _2354_ _2344_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4467_ _2306_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3418_ _1019_ _1024_ _1448_ _1083_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__o31a_1
X_4398_ _2186_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_37_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3349_ GCDdpath0.B_reg\[115\] _1325_ _1327_ _1385_ _1387_ VGND VGND VPWR VPWR _1388_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_70_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5019_ clknet_leaf_10_clk _0351_ _0095_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_55_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2720_ net328 GCDdpath0.B_reg\[46\] VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2651_ _0643_ _0701_ _0644_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2582_ _0608_ _0622_ _0628_ _0631_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__o32a_1
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4321_ net373 _2203_ _2201_ VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4252_ net268 _2154_ _2144_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3203_ _1089_ _1253_ _1032_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4183_ _2106_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3134_ _0746_ _0749_ _1183_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__o31a_1
XFILLER_0_145_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3065_ _1111_ _1112_ _1115_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3967_ net53 _1921_ _1898_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2918_ _0967_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
X_3898_ _1862_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2849_ GCDdpath0.B_reg\[83\] net369 VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4519_ GCDdpath0.B_reg\[28\] net177 _2342_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4870_ _2453_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3821_ _1794_ _1795_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3752_ _1736_ _1726_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2703_ net335 GCDdpath0.B_reg\[52\] VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__and2b_1
XFILLER_0_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3683_ _1677_ _0960_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2634_ _0680_ _0675_ _0678_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__or3b_1
XFILLER_0_3_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2565_ net291 GCDdpath0.B_reg\[12\] VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput268 net268 VGND VGND VPWR VPWR result_bits_data[107] sky130_fd_sc_hd__clkbuf_4
X_4304_ net379 _2191_ _2187_ VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__mux2_1
Xoutput279 net279 VGND VGND VPWR VPWR result_bits_data[117] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2496_ GCDdpath0.B_reg\[115\] GCDdpath0.B_reg\[114\] GCDdpath0.B_reg\[113\] GCDdpath0.B_reg\[112\]
+ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__or4_1
X_4235_ GCDdpath0.B_reg\[112\] net143 _2142_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4166_ net62 _2092_ _1287_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3117_ _0644_ _0653_ _0703_ _0643_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__a211o_1
X_4097_ GCDdpath0.B_reg\[13\] _2033_ _1834_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__mux2_1
X_3048_ GCDdpath0.B_reg\[117\] net279 VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4999_ clknet_leaf_21_clk _0331_ _0075_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4020_ net393 _0691_ _1966_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4922_ _2409_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4853_ _2451_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3804_ net78 _1781_ _1718_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4784_ _2439_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3735_ _0684_ _0708_ _0806_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3666_ _0922_ _1662_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__xnor2_1
X_2617_ net300 GCDdpath0.B_reg\[20\] VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3597_ _0906_ _1574_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__nor2_1
X_2548_ _0578_ _0585_ _0586_ _0587_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a311o_1
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2479_ _0523_ _0524_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or3_1
X_4218_ GCDdpath0.B_reg\[117\] net148 _2127_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4149_ _2078_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3520_ net122 _1432_ _1479_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3451_ GCDdpath0.B_reg\[103\] _1417_ _1418_ _1477_ _1387_ VGND VGND VPWR VPWR _1478_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3382_ _1284_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5121_ clknet_leaf_22_clk _0453_ _0197_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_88_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5052_ clknet_leaf_2_clk _0384_ _0128_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4003_ _0701_ _1938_ _0645_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4905_ _2459_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4836_ _2448_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4767_ _2437_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3718_ net91 _1707_ _1665_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4698_ _2425_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3649_ GCDdpath0.B_reg\[76\] _1648_ _1598_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 net210 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2951_ _0855_ _0859_ _1001_ _0850_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__o31a_1
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2882_ net364 GCDdpath0.B_reg\[79\] VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_40_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4621_ net258 net388 _2412_ net397 _2413_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ GCDdpath0.B_reg\[18\] net166 _2356_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3503_ net124 _1522_ _1468_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__mux2_1
X_4483_ GCDdpath0.B_reg\[39\] net189 _2314_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3434_ net266 _1462_ _1393_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3365_ net16 _1401_ _1337_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ clknet_leaf_29_clk _0436_ _0180_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3296_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__clkbuf_2
X_5035_ clknet_leaf_3_clk _0367_ _0111_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4819_ _2445_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput102 operands_bits_A[76] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
Xinput113 operands_bits_A[86] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
Xinput124 operands_bits_A[96] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput135 operands_bits_B[105] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
XFILLER_0_76_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput146 operands_bits_B[115] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_1
Xinput157 operands_bits_B[125] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
Xinput168 operands_bits_B[1] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
Xinput179 operands_bits_B[2] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_76_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3150_ _0795_ _0798_ _0799_ _1200_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3081_ GCDdpath0.B_reg\[122\] net285 VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_50_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3983_ _1764_ _1917_ _1933_ _1934_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2934_ _0963_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2865_ net359 GCDdpath0.B_reg\[74\] VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4604_ GCDdpath0.B_reg\[2\] net179 _1495_ VGND VGND VPWR VPWR _2402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ _0723_ _0720_ _0719_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4535_ GCDdpath0.B_reg\[23\] net172 _2342_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4466_ net326 _2305_ _2301_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3417_ _1084_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4397_ GCDdpath0.B_reg\[64\] net217 _2256_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3348_ _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3279_ _1299_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5018_ clknet_leaf_10_clk _0350_ _0094_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2650_ GCDdpath0.B_reg\[24\] net304 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2581_ _0629_ GCDdpath0.B_reg\[11\] VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4320_ GCDdpath0.B_reg\[87\] net242 _2199_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4251_ GCDdpath0.B_reg\[107\] net137 _2142_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3202_ _1038_ GCDdpath0.B_reg\[108\] _1037_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_52_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4182_ net394 _2105_ _1292_ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3133_ _0731_ _0745_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3064_ _1113_ _1114_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3966_ GCDdpath0.B_reg\[31\] _1920_ _1892_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2917_ net353 _0966_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3897_ _1860_ _1861_ _1609_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2848_ net369 GCDdpath0.B_reg\[83\] VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2779_ GCDdpath0.B_reg\[47\] net329 VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4518_ _2313_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4449_ net331 _2293_ _2287_ VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3820_ _0739_ _1772_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3751_ _0838_ _1186_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2702_ GCDdpath0.B_reg\[53\] net336 VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3682_ _0968_ _0972_ _1676_ _0967_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2633_ _0624_ _0638_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2564_ GCDdpath0.B_reg\[12\] net291 VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4303_ GCDdpath0.B_reg\[92\] net248 _2184_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__mux2_1
Xoutput269 net269 VGND VGND VPWR VPWR result_bits_data[108] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2495_ GCDdpath0.B_reg\[127\] GCDdpath0.B_reg\[126\] GCDdpath0.B_reg\[125\] GCDdpath0.B_reg\[124\]
+ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4234_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4165_ GCDdpath0.B_reg\[3\] _2091_ _1989_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3116_ _1163_ _1165_ _1166_ _0663_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4096_ _0618_ _2032_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_69_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3047_ _1093_ _1094_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__or3_2
XFILLER_0_78_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4998_ clknet_2_3__leaf_clk _0330_ _0074_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3949_ _1903_ _1905_ _1609_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_92_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4921_ _2461_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4852_ _2451_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3803_ GCDdpath0.B_reg\[54\] _1780_ _1684_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4783_ _2439_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3734_ _0719_ _0723_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__and2b_1
XFILLER_0_166_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3665_ _0987_ _1628_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2616_ _0665_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3596_ _1603_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2547_ _0591_ _0594_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2478_ _0525_ _0527_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or3_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4217_ _2130_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4148_ net354 _2077_ _2041_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4079_ _0617_ _2017_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3450_ _1471_ _1476_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3381_ net274 _1408_ _1413_ _1416_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5120_ clknet_leaf_14_clk _0452_ _0196_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5051_ clknet_leaf_1_clk _0383_ _0127_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4002_ _0645_ _0701_ _1938_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_148_Left_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4904_ _2459_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4835_ _2448_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4766_ _2437_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3717_ GCDdpath0.B_reg\[66\] _1706_ _1684_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4697_ _2425_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_157_Left_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3648_ _0929_ _1647_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3579_ net113 _1583_ _1479_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__o21a_1
XFILLER_0_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Left_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2950_ _0857_ _0860_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2881_ GCDdpath0.B_reg\[79\] net364 VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4620_ _2408_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__buf_2
XFILLER_0_84_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4551_ _2365_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_160_Right_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3502_ _1280_ _1498_ _1519_ _1521_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4482_ _2317_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3433_ net7 _1461_ _1337_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3364_ GCDdpath0.B_reg\[113\] _1395_ _1397_ _1400_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_55_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ clknet_leaf_29_clk _0435_ _0179_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _1287_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__clkbuf_4
X_5034_ clknet_leaf_6_clk _0366_ _0110_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4818_ _2445_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4749_ _2434_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput103 operands_bits_A[77] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
Xinput114 operands_bits_A[87] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
Xinput125 operands_bits_A[97] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
Xinput136 operands_bits_B[106] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_1
Xinput147 operands_bits_B[116] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_1
Xinput158 operands_bits_B[126] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput169 operands_bits_B[20] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_171_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3080_ net285 GCDdpath0.B_reg\[122\] VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3982_ GCDdpath0.B_reg\[28\] _1520_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2933_ _0967_ _0972_ _0983_ _0968_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2864_ _0913_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4603_ _2401_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2795_ _0759_ _0837_ _0845_ _0724_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_96_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4534_ _2353_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4465_ GCDdpath0.B_reg\[44\] net195 _2299_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3416_ _1027_ _1422_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4396_ _2227_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__buf_2
X_3347_ _1287_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__buf_2
X_3278_ _1284_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5017_ clknet_leaf_11_clk _0349_ _0093_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2580_ _0629_ GCDdpath0.B_reg\[11\] _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_112_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4250_ _2153_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__clkbuf_1
X_3201_ _1017_ _1019_ _1251_ _1040_ _1086_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_52_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4181_ net1 _2104_ _1287_ VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3132_ _0752_ _0754_ _1182_ _0813_ _0809_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__o311a_1
X_3063_ net274 GCDdpath0.B_reg\[112\] VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3965_ _1913_ _1919_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__xor2_1
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2916_ net353 _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3896_ net323 net64 _1615_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2847_ _0896_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2778_ _0773_ _0776_ _0777_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4517_ _2341_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4448_ GCDdpath0.B_reg\[49\] net200 _2285_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4379_ net355 _2243_ _2244_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3750_ net346 _1440_ _1733_ _1559_ _1735_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2701_ net336 GCDdpath0.B_reg\[53\] VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3681_ _0978_ _1675_ _0970_ _0972_ _0944_ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_171_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2632_ _0663_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2563_ _0610_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4302_ _2190_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput259 net259 VGND VGND VPWR VPWR operands_rdy sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2494_ GCDdpath0.B_reg\[123\] GCDdpath0.B_reg\[122\] GCDdpath0.B_reg\[121\] GCDdpath0.B_reg\[120\]
+ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or4_1
X_4233_ _1404_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4164_ _1175_ _2090_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3115_ net393 _0691_ _0665_ _0666_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__o31a_1
X_4095_ _0615_ _2018_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__nor2_1
X_3046_ _1095_ _1096_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4997_ clknet_leaf_21_clk _0329_ _0073_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3948_ net314 net55 _1904_ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3879_ net326 _1407_ _1846_ _1303_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _2461_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4851_ _2447_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ _0750_ _1775_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4782_ _2439_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3733_ _1720_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_635 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3664_ _1661_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2615_ net303 GCDdpath0.B_reg\[23\] VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3595_ net370 _1600_ _1602_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2546_ _0595_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nand2_1
X_2477_ GCDdpath0.B_reg\[35\] GCDdpath0.B_reg\[34\] GCDdpath0.B_reg\[33\] GCDdpath0.B_reg\[32\]
+ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4216_ net280 _2128_ _2129_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4147_ net95 _2076_ _2029_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4078_ _0631_ _2016_ _0632_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ _1055_ GCDdpath0.B_reg\[103\] _1061_ _1078_ _1079_ VGND VGND VPWR VPWR _1080_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_84_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_174_Right_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3380_ net15 _1414_ _1415_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5050_ clknet_leaf_1_clk _0382_ _0126_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4001_ net305 net46 _1406_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4903_ _2459_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4834_ _2448_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4765_ _2433_ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__buf_2
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3716_ _0949_ _1705_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4696_ _2425_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3647_ _0991_ _1629_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3578_ GCDdpath0.B_reg\[86\] _1296_ _1587_ _1303_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2529_ GCDdpath0.B_reg\[0\] VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__inv_2
X_5179_ clknet_leaf_1_clk _0511_ _0255_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2880_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4550_ net298 _2364_ _2358_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3501_ GCDdpath0.B_reg\[96\] _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__and2_1
X_4481_ net322 _2315_ _2316_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3432_ _1459_ _1460_ _1395_ GCDdpath0.B_reg\[105\] VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3363_ _1398_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5102_ clknet_leaf_38_clk _0434_ _0178_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_55_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _1339_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_1
X_5033_ clknet_leaf_8_clk _0365_ _0109_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4817_ _2445_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4748_ _2434_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_151_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4679_ _2419_ VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput104 operands_bits_A[78] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
Xinput115 operands_bits_A[88] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xinput126 operands_bits_A[98] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xinput137 operands_bits_B[107] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xinput148 operands_bits_B[117] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput159 operands_bits_B[127] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3981_ _0658_ _0705_ _1916_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__nand3_1
XFILLER_0_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2932_ _0979_ _0982_ _0969_ _0973_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_42_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2863_ net360 GCDdpath0.B_reg\[75\] VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4602_ net321 _2400_ _2044_ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2794_ _0726_ _0838_ _0730_ _0844_ _0728_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_96_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4533_ net304 _2352_ _2344_ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ _2304_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3415_ _1017_ _1018_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4395_ _2255_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3346_ _1382_ _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3277_ _1293_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_29_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ clknet_leaf_17_clk _0348_ _0092_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_15_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3200_ _1250_ _1026_ _1020_ _1023_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4180_ GCDdpath0.B_reg\[0\] _2103_ _1279_ VGND VGND VPWR VPWR _2104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3131_ _0742_ _1181_ _0755_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_173_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3062_ GCDdpath0.B_reg\[112\] net274 VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3964_ _0649_ _0660_ _1918_ _0698_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2915_ GCDdpath0.B_reg\[69\] VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3895_ GCDdpath0.B_reg\[41\] _1859_ _1620_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2846_ net366 _0895_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2777_ net329 GCDdpath0.B_reg\[47\] VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4516_ net309 _2340_ _2330_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4447_ _2292_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4378_ _2186_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__buf_2
X_3329_ net280 _1324_ _1368_ _1370_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_146_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2700_ _0747_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3680_ _0981_ _1674_ _0950_ _0951_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2631_ _0672_ _0675_ _0678_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2562_ _0611_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4301_ net380 _2189_ _2187_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2493_ GCDdpath0.B_reg\[119\] GCDdpath0.B_reg\[118\] GCDdpath0.B_reg\[117\] GCDdpath0.B_reg\[116\]
+ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__or4_1
X_4232_ _2140_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_4_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_4163_ _0578_ _0585_ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3114_ _0664_ _0667_ _0670_ _1164_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__or4_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4094_ _2031_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__clkbuf_1
X_3045_ GCDdpath0.B_reg\[114\] net276 VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_69_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4996_ clknet_leaf_24_clk _0328_ _0072_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3947_ _1405_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_82_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3878_ _1843_ _1437_ _1620_ _1845_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2829_ net371 GCDdpath0.B_reg\[85\] VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _2450_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3801_ net338 _1349_ _1778_ _1779_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_64_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4781_ _2439_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3732_ net348 _1719_ _1687_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3663_ net359 _1660_ _1602_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2614_ GCDdpath0.B_reg\[23\] net303 VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__and2b_1
X_3594_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2545_ net332 GCDdpath0.B_reg\[4\] VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2476_ GCDdpath0.B_reg\[47\] _0526_ GCDdpath0.B_reg\[45\] GCDdpath0.B_reg\[44\] VGND
+ VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4215_ _2082_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4146_ _1764_ _2068_ _2074_ _2075_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4077_ _0621_ _2015_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3028_ _1057_ _1058_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4979_ clknet_leaf_27_clk _0311_ _0055_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4000_ net306 _1408_ _1948_ _1949_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4902_ _2459_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4833_ _2448_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4764_ _2436_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3715_ _0981_ _1674_ _0951_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4695_ _2425_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3646_ net362 _1440_ _1645_ _1559_ _1646_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3577_ _1579_ _1586_ _1300_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2528_ GCDdpath0.B_reg\[1\] net299 VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5178_ clknet_leaf_3_clk _0510_ _0254_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4129_ _1764_ _2014_ _2059_ _2060_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3500_ _1398_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4480_ _2272_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__buf_2
X_3431_ _1250_ _1448_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3362_ _1111_ _1112_ _1113_ _1396_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5101_ clknet_leaf_38_clk _0433_ _0177_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_55_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ net285 _1338_ _1322_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5032_ clknet_leaf_8_clk _0364_ _0108_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4816_ _2445_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4747_ _2434_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4678_ _2422_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3629_ _0925_ _0936_ _1631_ _0935_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput105 operands_bits_A[79] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xinput116 operands_bits_A[89] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xinput127 operands_bits_A[99] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput138 operands_bits_B[108] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
Xinput149 operands_bits_B[118] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_158_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3980_ _1932_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2931_ _0978_ _0980_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2862_ GCDdpath0.B_reg\[75\] net360 VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4601_ GCDdpath0.B_reg\[3\] net190 _1495_ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2793_ _0711_ _0715_ _0839_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_96_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4532_ GCDdpath0.B_reg\[24\] net173 _2342_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4463_ net327 _2303_ _2301_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3414_ _1293_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4394_ net349 _2254_ _2244_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3345_ _1095_ _1383_ _1121_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__a21oi_1
X_3276_ _1323_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5015_ clknet_leaf_16_clk _0347_ _0091_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_153_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_169_Right_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3130_ _0734_ _0736_ _0744_ _1180_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_59_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3061_ net275 GCDdpath0.B_reg\[113\] VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3963_ _0700_ _1917_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__or2b_1
XFILLER_0_86_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2914_ _0960_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3894_ _0788_ _1858_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__xor2_1
XFILLER_0_169_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2845_ net366 _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2776_ net328 VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4515_ GCDdpath0.B_reg\[29\] net178 _2328_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4446_ net333 _2291_ _2287_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4377_ GCDdpath0.B_reg\[70\] net224 _2242_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3328_ net21 _1305_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_146_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _0572_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_107_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2630_ _0679_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2561_ net376 GCDdpath0.B_reg\[8\] VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4300_ GCDdpath0.B_reg\[93\] net249 _2184_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2492_ _0530_ _0531_ _0535_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4231_ net275 _2139_ _2129_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__mux2_1
X_4162_ _2089_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_1
X_3113_ _0693_ _0536_ _0669_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4093_ net293 _2030_ _1992_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__mux2_1
X_3044_ net276 GCDdpath0.B_reg\[114\] VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_69_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4995_ clknet_leaf_21_clk _0327_ _0071_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3946_ GCDdpath0.B_reg\[33\] _1902_ _1834_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3877_ _1825_ _1844_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2828_ _0862_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2759_ _0739_ _0743_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4429_ net338 _2279_ _2273_ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ net79 _1583_ _1517_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4780_ _2439_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3731_ net89 _1717_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_172_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3662_ net100 _1659_ _1565_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2613_ net393 GCDdpath0.B_reg\[22\] VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__xor2_2
XFILLER_0_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3593_ _1291_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2544_ GCDdpath0.B_reg\[4\] net332 VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or2b_1
XFILLER_0_140_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2475_ GCDdpath0.B_reg\[46\] VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_103_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4214_ GCDdpath0.B_reg\[118\] net149 _2127_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4145_ GCDdpath0.B_reg\[6\] _1398_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_3_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4076_ _0628_ _2014_ _0608_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3027_ _1068_ _1076_ _1077_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4978_ clknet_leaf_29_clk _0310_ _0054_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3929_ _0765_ _1821_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4901_ _2454_ VGND VGND VPWR VPWR _2459_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4832_ _2448_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4763_ _2436_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3714_ _1704_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4694_ _2425_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3645_ net103 _1506_ _1355_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3576_ _0889_ _1585_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2527_ GCDdpath0.B_reg\[2\] net310 VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_114_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5177_ clknet_leaf_3_clk _0509_ _0253_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4128_ GCDdpath0.B_reg\[8\] _1398_ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4059_ net296 GCDdpath0.B_reg\[17\] VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3430_ _1299_ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3361_ _1298_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5100_ clknet_leaf_28_clk _0432_ _0176_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dfrtp_4
X_3292_ net26 _1335_ _1337_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ clknet_leaf_8_clk _0363_ _0107_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4815_ _2440_ VGND VGND VPWR VPWR _2445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4746_ _2434_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4677_ _2422_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_151_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3628_ _0994_ _0927_ _1630_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3559_ net115 _1570_ _1565_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput106 operands_bits_A[7] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xinput117 operands_bits_A[8] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput128 operands_bits_A[9] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput139 operands_bits_B[109] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2930_ _0952_ _0954_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__and2b_1
XFILLER_0_168_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2861_ _0879_ _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__or2_2
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4600_ _2399_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2792_ net392 _0840_ _0841_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4531_ _2351_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4462_ GCDdpath0.B_reg\[45\] net196 _2299_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3413_ net269 _1440_ _1443_ _1354_ _1444_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4393_ GCDdpath0.B_reg\[65\] net218 _2242_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3344_ _1120_ _1358_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3275_ net287 _1321_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5014_ clknet_leaf_11_clk _0346_ _0090_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4729_ _2426_ VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3060_ GCDdpath0.B_reg\[113\] net275 VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3962_ _0705_ _1916_ _0658_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2913_ _0962_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3893_ _0791_ _1823_ _0790_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2844_ GCDdpath0.B_reg\[80\] VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2775_ _0781_ _0824_ _0825_ _0779_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4514_ _2339_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4445_ GCDdpath0.B_reg\[50\] net202 _2285_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4376_ _2227_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__buf_2
X_3327_ _0572_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ net289 _1294_ _1304_ _1307_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_163_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _0855_ _0860_ _1238_ _1239_ net381 VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_124_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2560_ GCDdpath0.B_reg\[8\] net376 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2491_ _0537_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or2_1
X_4230_ GCDdpath0.B_reg\[113\] net144 _2127_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__mux2_1
X_4161_ net332 _2088_ _2041_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__mux2_1
X_3112_ _1160_ _1162_ _0672_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__a21o_1
X_4092_ net34 _2028_ _2029_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3043_ net277 GCDdpath0.B_reg\[115\] VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4994_ clknet_leaf_22_clk _0326_ _0070_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3945_ _0768_ _1901_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_82_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3876_ _0775_ _1824_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2827_ _0870_ _0874_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__or3_1
XFILLER_0_171_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2758_ GCDdpath0.B_reg\[54\] net337 VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2689_ net333 GCDdpath0.B_reg\[50\] VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_148_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4428_ GCDdpath0.B_reg\[55\] net207 _2270_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4359_ net361 _2229_ _2230_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3730_ _1336_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3661_ GCDdpath0.B_reg\[74\] _1658_ _1598_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2612_ _0646_ _0652_ _0655_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__or4_2
X_3592_ net111 _1599_ _1565_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ _0592_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2474_ GCDdpath0.B_reg\[43\] GCDdpath0.B_reg\[42\] GCDdpath0.B_reg\[41\] GCDdpath0.B_reg\[40\]
+ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or4_1
XFILLER_0_55_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4213_ _1405_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__buf_2
XFILLER_0_103_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4144_ _0590_ _2067_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4075_ _0613_ _2013_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3026_ _1062_ _1066_ _1065_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_84_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4977_ clknet_leaf_29_clk _0309_ _0053_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3928_ _1887_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3859_ GCDdpath0.B_reg\[47\] _1325_ _1409_ _1829_ _1415_ VGND VGND VPWR VPWR _1830_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4900_ _2458_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4831_ _2448_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4762_ _2436_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3713_ net351 _1703_ _1687_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4693_ _2419_ VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3644_ GCDdpath0.B_reg\[77\] _1644_ _1442_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3575_ _0885_ _1577_ _1578_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2526_ GCDdpath0.B_reg\[125\] net288 VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_114_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5176_ clknet_leaf_3_clk _0508_ _0252_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dfrtp_4
X_4127_ _0613_ _2013_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4058_ _1999_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3009_ _1058_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3360_ _1111_ _1112_ _1113_ _1396_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__nor4_1
XFILLER_0_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__clkbuf_4
X_5030_ clknet_leaf_7_clk _0362_ _0106_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_45_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4814_ _2444_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4745_ _2434_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4676_ _2422_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3627_ _0991_ _1629_ _0929_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3558_ GCDdpath0.B_reg\[88\] _1569_ _1482_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2509_ GCDdpath0.B_reg\[95\] GCDdpath0.B_reg\[94\] GCDdpath0.B_reg\[93\] GCDdpath0.B_reg\[92\]
+ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__or4_1
X_3489_ net384 net125 _1496_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__mux2_1
Xinput107 operands_bits_A[80] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput118 operands_bits_A[90] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_1
Xinput129 operands_bits_B[0] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_5159_ clknet_leaf_8_clk _0491_ _0235_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2860_ _0894_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2791_ GCDdpath0.B_reg\[59\] net342 VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Left_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4530_ net305 _2350_ _2344_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4461_ _2302_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3412_ net10 _1288_ _1355_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4392_ _2253_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3343_ _1093_ _1094_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3274_ _1292_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_163_Left_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5013_ clknet_leaf_11_clk _0345_ _0089_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_165_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_172_Left_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2989_ _1038_ GCDdpath0.B_reg\[108\] VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__or2_2
XFILLER_0_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4728_ _2430_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4659_ _2420_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3961_ _0646_ _0655_ _1915_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__or3_1
XFILLER_0_159_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2912_ net356 _0961_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3892_ _1857_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2843_ _0880_ _0881_ _0885_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2774_ _0780_ _0784_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4513_ net311 _2338_ _2330_ VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4444_ _2290_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4375_ _2241_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3326_ GCDdpath0.B_reg\[118\] _1325_ _1327_ _1367_ _1303_ VGND VGND VPWR VPWR _1368_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_146_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ net30 _1305_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3188_ GCDdpath0.B_reg\[94\] _0850_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2490_ _0538_ _0539_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4160_ net73 _2087_ _2029_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__mux2_1
X_3111_ _0675_ _1161_ _0687_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__o21a_1
X_4091_ _1286_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__buf_2
XFILLER_0_171_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3042_ GCDdpath0.B_reg\[115\] net277 VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__nor2b_1
XTAP_TAPCELL_ROW_19_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4993_ clknet_leaf_22_clk _0325_ _0069_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3944_ _0763_ _1888_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3875_ GCDdpath0.B_reg\[44\] VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2826_ _0875_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2757_ _0684_ _0708_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a21o_2
XFILLER_0_143_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2688_ GCDdpath0.B_reg\[50\] net333 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_148_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4427_ _2278_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _2186_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__buf_2
X_3309_ _0571_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ net383 _2180_ _2172_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3660_ _0918_ _1657_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2611_ _0658_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or2b_1
XFILLER_0_153_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3591_ GCDdpath0.B_reg\[84\] _1597_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ net343 GCDdpath0.B_reg\[5\] VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2473_ GCDdpath0.B_reg\[39\] GCDdpath0.B_reg\[38\] GCDdpath0.B_reg\[37\] GCDdpath0.B_reg\[36\]
+ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4212_ _2126_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4143_ _2073_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4074_ _0599_ _0601_ _0604_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_104_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3025_ _1072_ _0553_ _1073_ _1045_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__o311a_1
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4976_ clknet_leaf_29_clk _0308_ _0052_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_164_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3927_ net317 _1886_ _1841_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3858_ _0770_ _1828_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2809_ GCDdpath0.B_reg\[93\] net380 VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3789_ net339 _1768_ _1745_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4830_ _2447_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4761_ _2436_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3712_ net92 _1702_ _1665_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4692_ _2424_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3643_ _0926_ _1643_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3574_ net373 _1445_ _1582_ _1584_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2525_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5175_ clknet_leaf_13_clk _0507_ _0251_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dfrtp_4
X_4126_ _1509_ _2054_ _2057_ _2058_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o22a_1
X_4057_ net297 _1998_ _1992_ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3008_ net263 GCDdpath0.B_reg\[102\] VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4959_ clknet_leaf_34_clk _0291_ _0035_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_49_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput380 net380 VGND VGND VPWR VPWR result_bits_data[93] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_674 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_164_Right_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3290_ _1286_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4813_ _2444_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4744_ _2433_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4675_ _2422_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3626_ _0923_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3557_ _1551_ _1568_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2508_ GCDdpath0.B_reg\[91\] GCDdpath0.B_reg\[90\] GCDdpath0.B_reg\[89\] GCDdpath0.B_reg\[88\]
+ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__or4_1
XFILLER_0_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3488_ _1508_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__clkbuf_4
Xinput108 operands_bits_A[81] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
Xinput119 operands_bits_A[91] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlymetal6s2s_1
X_5158_ clknet_leaf_7_clk _0490_ _0234_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dfrtp_4
X_4109_ _1281_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__buf_2
X_5089_ clknet_leaf_34_clk _0421_ _0165_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2790_ net342 GCDdpath0.B_reg\[59\] VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4460_ net328 _2300_ _2301_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3411_ GCDdpath0.B_reg\[108\] _1441_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4391_ net350 _2252_ _2244_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3342_ _1381_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3273_ net28 _1320_ _1302_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5012_ clknet_leaf_16_clk _0344_ _0088_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2988_ _1038_ GCDdpath0.B_reg\[108\] VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4727_ _2430_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4658_ _2419_ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 operands_bits_A[65] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
X_3609_ net368 _1294_ _1614_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4589_ GCDdpath0.B_reg\[7\] net234 _2384_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3960_ _0690_ _0692_ _0695_ _1914_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2911_ net356 _0961_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__nor2_1
X_3891_ net324 _1856_ _1841_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2842_ _0889_ _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2773_ _0787_ _0790_ _0782_ _0785_ _0786_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_170_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4512_ GCDdpath0.B_reg\[30\] net180 _2328_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4443_ net334 _2289_ _2287_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4374_ net356 _2240_ _2230_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3325_ _1361_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__nor2_1
X_3256_ _0572_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_146_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _0856_ _0859_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap390 _1177_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3110_ _0677_ _0681_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nand2_1
X_4090_ _1464_ _2019_ _2026_ _2027_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3041_ _1043_ _1080_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4992_ clknet_leaf_24_clk _0324_ _0068_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3943_ _1900_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3874_ _1842_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2825_ _0872_ GCDdpath0.B_reg\[88\] VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2756_ _0759_ _0806_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__or2_2
XFILLER_0_171_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2687_ _0734_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_148_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4426_ net339 _2277_ _2273_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_165_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ GCDdpath0.B_reg\[76\] net230 _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__mux2_1
X_3308_ GCDdpath0.B_reg\[120\] _1351_ _1296_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ GCDdpath0.B_reg\[96\] net252 _2170_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _1159_ _1282_ _1283_ _1289_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2610_ _0659_ _0660_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and2b_1
X_3590_ _1318_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2541_ GCDdpath0.B_reg\[5\] net343 VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2b_1
XFILLER_0_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2472_ _0519_ _0520_ _0521_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4211_ net281 _2125_ _2115_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4142_ _2071_ _2072_ _1609_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4073_ GCDdpath0.B_reg\[14\] VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3024_ _1048_ _1049_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_104_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4975_ clknet_leaf_29_clk _0307_ _0051_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3926_ net58 _1885_ _1817_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3857_ _1208_ _0777_ _1826_ _1827_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2808_ net380 GCDdpath0.B_reg\[93\] VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3788_ net80 _1767_ _1718_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2739_ GCDdpath0.B_reg\[40\] net322 VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4409_ _2265_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4760_ _2436_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3711_ _0564_ _1701_ _1684_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4691_ _2424_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3642_ _1636_ _1630_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3573_ net114 _1583_ _1479_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2524_ GCDdpath0.B_reg\[126\] net289 VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5174_ clknet_leaf_13_clk _0506_ _0250_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dfrtp_4
X_4125_ net399 _1516_ _1353_ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__a21o_1
X_4056_ net38 _1997_ _1984_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3007_ GCDdpath0.B_reg\[102\] net263 VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4958_ clknet_leaf_34_clk _0290_ _0034_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3909_ _0795_ _1871_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_173_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4889_ _2457_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput370 net370 VGND VGND VPWR VPWR result_bits_data[84] sky130_fd_sc_hd__clkbuf_4
Xoutput381 net381 VGND VGND VPWR VPWR result_bits_data[94] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4812_ _2444_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4743_ _2408_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__buf_2
XFILLER_0_127_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4674_ _2422_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3625_ _0986_ _1627_ _0941_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3556_ _1550_ _1012_ _1527_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2507_ GCDdpath0.B_reg\[83\] GCDdpath0.B_reg\[82\] GCDdpath0.B_reg\[81\] GCDdpath0.B_reg\[80\]
+ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or4_1
X_3487_ _1386_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__buf_2
Xinput109 operands_bits_A[82] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_5157_ clknet_leaf_8_clk _0489_ _0233_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dfrtp_4
X_4108_ net282 net23 _1406_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__mux2_1
X_5088_ clknet_leaf_36_clk _0420_ _0164_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dfrtp_4
X_4039_ _0536_ _1982_ _1892_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_167_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3410_ _1295_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__buf_4
X_4390_ GCDdpath0.B_reg\[66\] net219 _2242_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3341_ net278 _1380_ _1322_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__mux2_1
X_3272_ GCDdpath0.B_reg\[124\] _1317_ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__mux2_1
X_5011_ clknet_leaf_16_clk _0343_ _0087_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2987_ net269 VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4726_ _2430_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4657_ _2408_ VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_131_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput80 operands_bits_A[56] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3608_ net109 _1609_ _1612_ _1613_ _1407_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput91 operands_bits_A[66] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
X_4588_ _2391_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3539_ _0865_ _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2910_ GCDdpath0.B_reg\[71\] VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3890_ net65 _1855_ _1817_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2841_ _0890_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2772_ _0818_ _0822_ _0779_ _0792_ _0805_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4511_ _2337_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4442_ GCDdpath0.B_reg\[51\] net203 _2285_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4373_ GCDdpath0.B_reg\[71\] net225 _2228_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3324_ _1109_ _1125_ _1360_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3255_ _0516_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _1234_ _1235_ _1236_ _0862_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4709_ _2428_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap391 _0758_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3040_ _1081_ _1030_ _1035_ _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_159_Right_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4991_ clknet_leaf_23_clk _0323_ _0067_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3942_ net315 _1899_ _1841_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3873_ net327 _1840_ _1841_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2824_ net375 GCDdpath0.B_reg\[89\] VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_30_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2755_ _0769_ _0779_ _0792_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or4_1
XFILLER_0_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2686_ _0735_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4425_ GCDdpath0.B_reg\[56\] net208 _2270_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4356_ _2227_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3307_ _1139_ _1350_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__xnor2_1
X_4287_ _2179_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_126_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ GCDdpath0.B_reg\[127\] _1285_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__o21ai_1
X_3169_ _0928_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_169_Left_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2540_ _0588_ _0589_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2471_ GCDdpath0.B_reg\[51\] GCDdpath0.B_reg\[50\] GCDdpath0.B_reg\[49\] GCDdpath0.B_reg\[48\]
+ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4210_ GCDdpath0.B_reg\[119\] net150 _2113_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__mux2_1
X_4141_ net365 net106 _1904_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4072_ _2011_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_160_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3023_ _1052_ _1050_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4974_ clknet_leaf_27_clk _0306_ _0050_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3925_ GCDdpath0.B_reg\[36\] _1884_ _1810_ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3856_ _0827_ _0526_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2807_ _0856_ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3787_ _1764_ _1747_ _1765_ _1766_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_119_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2738_ net322 GCDdpath0.B_reg\[40\] VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2669_ GCDdpath0.B_reg\[62\] net346 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4408_ net345 _2264_ _2258_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4339_ _2216_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3710_ _1699_ _1700_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__nand2_1
X_4690_ _2424_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3641_ _1642_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3572_ _0516_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2523_ net31 _0517_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5173_ clknet_leaf_4_clk _0505_ _0249_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dfrtp_4
X_4124_ _1511_ _2055_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__nor3_1
Xinput1 operands_bits_A[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_4055_ GCDdpath0.B_reg\[18\] _1996_ _1989_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
X_3006_ _1055_ GCDdpath0.B_reg\[103\] VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4957_ clknet_leaf_36_clk _0289_ _0033_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3908_ _0798_ _1870_ _0797_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_163_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4888_ _2457_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3839_ net72 _1811_ _1718_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput360 net360 VGND VGND VPWR VPWR result_bits_data[75] sky130_fd_sc_hd__clkbuf_4
Xoutput371 net371 VGND VGND VPWR VPWR result_bits_data[85] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput382 net382 VGND VGND VPWR VPWR result_bits_data[95] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_124_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4811_ _2444_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4742_ _2432_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4673_ _2422_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3624_ _0808_ _0848_ _0975_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3555_ _1567_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2506_ GCDdpath0.B_reg\[87\] GCDdpath0.B_reg\[86\] GCDdpath0.B_reg\[85\] GCDdpath0.B_reg\[84\]
+ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3486_ net385 _1440_ _1505_ _1354_ _1507_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__o221a_1
X_5156_ clknet_leaf_9_clk _0488_ _0232_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4107_ _2042_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__clkbuf_1
X_5087_ clknet_leaf_34_clk _0419_ _0163_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4038_ _0668_ _1964_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3340_ net19 _1379_ _1337_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3271_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__clkbuf_4
X_5010_ clknet_leaf_15_clk _0342_ _0086_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2986_ net270 GCDdpath0.B_reg\[109\] VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_146_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4725_ _2430_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4656_ _2418_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_141_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput70 operands_bits_A[47] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
X_3607_ GCDdpath0.B_reg\[82\] _1281_ _1386_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput81 operands_bits_A[57] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4587_ net376 _2390_ _2386_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput92 operands_bits_A[67] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3538_ _0867_ _1552_ _0868_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_168_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3469_ net2 _1492_ _1468_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5139_ clknet_leaf_15_clk _0471_ _0215_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_150_Left_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2840_ GCDdpath0.B_reg\[87\] net373 VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_14_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2771_ _0819_ _0820_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4510_ net312 _2336_ _2330_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4441_ _2288_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4372_ _2239_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3323_ _1357_ _1365_ _1294_ net281 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3254_ GCDdpath0.B_reg\[126\] _1296_ _1301_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_146_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3185_ _0864_ _0867_ _0863_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_163_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2969_ GCDdpath0.B_reg\[106\] net267 VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4708_ _2426_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4639_ _2416_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4990_ clknet_leaf_24_clk _0322_ _0066_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3941_ net56 _1897_ _1898_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3872_ _1601_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2823_ _0871_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2754_ _0795_ _0798_ _0801_ _0804_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2685_ GCDdpath0.B_reg\[49\] net331 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4424_ _2276_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4355_ _1404_ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_165_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _1118_ _1127_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4286_ net384 _2178_ _2172_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _1287_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168_ net356 _0961_ _1217_ _1218_ _0958_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3099_ _1141_ _1144_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2470_ GCDdpath0.B_reg\[55\] GCDdpath0.B_reg\[54\] GCDdpath0.B_reg\[53\] GCDdpath0.B_reg\[52\]
+ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__or4_1
XFILLER_0_167_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4140_ GCDdpath0.B_reg\[7\] _2070_ _1834_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4071_ net295 _2010_ _1992_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3022_ net386 GCDdpath0.B_reg\[99\] VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_160_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4973_ clknet_leaf_37_clk _0305_ _0049_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3924_ _1869_ _1883_ VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3855_ _0773_ _0776_ _1825_ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2806_ GCDdpath0.B_reg\[92\] net379 VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__and2b_1
XFILLER_0_61_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3786_ GCDdpath0.B_reg\[56\] _1520_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_119_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2737_ _0786_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2668_ GCDdpath0.B_reg\[63\] net347 VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4407_ GCDdpath0.B_reg\[61\] net214 _2256_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2599_ GCDdpath0.B_reg\[30\] net311 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4338_ net368 _2214_ _2215_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__mux2_1
X_4269_ net263 _2166_ _2158_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3640_ net363 _1641_ _1602_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3571_ GCDdpath0.B_reg\[87\] _1285_ _1549_ _1581_ _1536_ VGND VGND VPWR VPWR _1582_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2522_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5172_ clknet_leaf_4_clk _0504_ _0248_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dfrtp_4
X_4123_ _0611_ _2014_ _0610_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__a21oi_1
Xinput2 operands_bits_A[100] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_4054_ _1963_ _1995_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__and2b_1
X_3005_ _1055_ GCDdpath0.B_reg\[103\] VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4956_ clknet_leaf_35_clk _0288_ _0032_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3907_ _0833_ _1869_ _0800_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_138_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4887_ _2454_ VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_173_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3838_ GCDdpath0.B_reg\[49\] _1809_ _1810_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3769_ net342 _1539_ _1751_ _1306_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput350 net350 VGND VGND VPWR VPWR result_bits_data[66] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput361 net361 VGND VGND VPWR VPWR result_bits_data[76] sky130_fd_sc_hd__clkbuf_4
Xoutput372 net372 VGND VGND VPWR VPWR result_bits_data[86] sky130_fd_sc_hd__clkbuf_4
Xoutput383 net383 VGND VGND VPWR VPWR result_bits_data[96] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_27_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4810_ _2444_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4741_ _2432_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4672_ _2419_ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3623_ net366 _1408_ _1625_ _1626_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3554_ net375 _1566_ _1489_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2505_ _0549_ _0550_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or3_1
X_3485_ net126 _1506_ _1355_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__or3_1
X_5155_ clknet_leaf_9_clk _0487_ _0231_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4106_ net291 _2040_ _2041_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__mux2_1
X_5086_ clknet_leaf_34_clk _0418_ _0162_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4037_ _1509_ _1977_ _1980_ _1981_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4939_ clknet_leaf_45_clk _0271_ _0015_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_859 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3270_ _1278_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2985_ GCDdpath0.B_reg\[109\] net270 VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4724_ _2430_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4655_ _2418_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput60 operands_bits_A[38] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_82_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3606_ _1574_ _1611_ _1296_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput71 operands_bits_A[48] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4586_ GCDdpath0.B_reg\[8\] net245 _2384_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__mux2_1
Xinput82 operands_bits_A[58] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput93 operands_bits_A[68] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlymetal6s2s_1
X_3537_ _0874_ _1551_ _0875_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3468_ GCDdpath0.B_reg\[100\] _1491_ _1482_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__mux2_1
X_3399_ net13 _1432_ _1369_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_129_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5138_ clknet_leaf_13_clk _0470_ _0214_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5069_ clknet_leaf_45_clk _0401_ _0145_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_165_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_164_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2770_ net316 GCDdpath0.B_reg\[35\] VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or2b_1
XFILLER_0_143_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4440_ net335 _2286_ _2287_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4371_ net357 _2238_ _2230_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3322_ _1282_ _1362_ _1363_ _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3253_ _1302_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3184_ _0870_ _0871_ _0877_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_163_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2968_ net267 GCDdpath0.B_reg\[106\] VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__and2b_1
XFILLER_0_162_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4707_ _2427_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2899_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__inv_2
X_4638_ _2416_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4569_ GCDdpath0.B_reg\[13\] net161 _2370_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_173_Right_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput250 operands_bits_B[94] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3940_ _1286_ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3871_ net68 _1839_ _1817_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2822_ _0872_ GCDdpath0.B_reg\[88\] VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2753_ _0802_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2684_ GCDdpath0.B_reg\[48\] net330 VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4423_ net340 _2275_ _2273_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4354_ _2226_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_165_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _1322_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__buf_2
X_4285_ GCDdpath0.B_reg\[97\] net253 _2170_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _1286_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__clkbuf_2
X_3167_ _0959_ _0968_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3098_ _0577_ _1145_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4070_ net36 _2009_ _1984_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3021_ net385 VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4972_ clknet_leaf_27_clk _0304_ _0048_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3923_ _0804_ _1822_ VGND VGND VPWR VPWR _1883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3854_ _0775_ _1824_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2805_ net379 GCDdpath0.B_reg\[92\] VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3785_ _0714_ _1724_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2736_ GCDdpath0.B_reg\[41\] net323 VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2667_ _0711_ _0714_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__or3_1
X_4406_ _2263_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2598_ net311 GCDdpath0.B_reg\[30\] VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__or2b_1
X_4337_ _2186_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4268_ GCDdpath0.B_reg\[102\] net132 _2156_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3219_ _1267_ _1131_ _1269_ _1129_ _1149_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_2_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4199_ net286 _2117_ _2115_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_173_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3570_ _0892_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2521_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5171_ clknet_leaf_5_clk _0503_ _0247_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4122_ _0610_ _0611_ _2014_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ _0673_ _1994_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__nand2_1
Xinput3 operands_bits_A[101] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_0_127_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3004_ net264 VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4955_ clknet_leaf_35_clk _0287_ _0031_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3906_ _0804_ _1822_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4886_ _2456_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3837_ _1318_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3768_ _1750_ _1281_ _1437_ GCDdpath0.B_reg\[59\] VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2719_ net329 GCDdpath0.B_reg\[47\] VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3699_ net353 _1539_ _1691_ _1306_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput340 net340 VGND VGND VPWR VPWR result_bits_data[57] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput351 net351 VGND VGND VPWR VPWR result_bits_data[67] sky130_fd_sc_hd__buf_2
Xoutput362 net362 VGND VGND VPWR VPWR result_bits_data[77] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput373 net373 VGND VGND VPWR VPWR result_bits_data[87] sky130_fd_sc_hd__clkbuf_4
Xoutput384 net384 VGND VGND VPWR VPWR result_bits_data[97] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4740_ _2432_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4671_ _2421_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3622_ net107 _1414_ _1415_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3553_ net116 _1564_ _1565_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2504_ _0551_ _0552_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__or3_1
X_3484_ _1302_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5154_ clknet_leaf_12_clk _0486_ _0230_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4105_ _1291_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__buf_2
X_5085_ clknet_leaf_36_clk _0417_ _0161_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4036_ GCDdpath0.B_reg\[21\] _1516_ _1353_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4938_ clknet_leaf_43_clk _0270_ _0014_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4869_ _2453_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2984_ _1029_ _1030_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4723_ _2430_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_170_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4654_ _2418_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput50 operands_bits_A[29] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
X_3605_ _0909_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput61 operands_bits_A[39] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
X_4585_ _2389_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
Xinput72 operands_bits_A[49] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XFILLER_0_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput83 operands_bits_A[59] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xinput94 operands_bits_A[69] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3536_ _1012_ _1527_ _1550_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_168_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3467_ _1064_ _1473_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3398_ _0516_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__clkbuf_2
X_5137_ clknet_leaf_25_clk _0469_ _0213_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dfrtp_4
X_5068_ clknet_leaf_46_clk _0400_ _0144_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4019_ _0694_ _1965_ _0664_ _0669_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4370_ GCDdpath0.B_reg\[72\] net226 _2228_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3321_ GCDdpath0.B_reg\[119\] _1313_ _1288_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3252_ _1287_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3183_ _1232_ _1233_ _0878_ _0891_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2967_ GCDdpath0.B_reg\[107\] net268 VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4706_ _2427_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2898_ _0947_ _0948_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__nor2_1
X_4637_ _2416_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4568_ _2377_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3519_ GCDdpath0.B_reg\[94\] _1417_ _1418_ _1535_ _1536_ VGND VGND VPWR VPWR _1537_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4499_ GCDdpath0.B_reg\[34\] net184 _2328_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput240 operands_bits_B[85] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 operands_bits_B[95] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_106_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ GCDdpath0.B_reg\[45\] _1838_ _1810_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2821_ net374 VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2752_ net317 GCDdpath0.B_reg\[36\] VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2683_ _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4422_ GCDdpath0.B_reg\[57\] net209 _2270_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4353_ net362 _2225_ _2215_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ net25 _1341_ _1342_ _1348_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_165_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4284_ _2177_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_129_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3235_ _0518_ _0569_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_126_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3166_ net353 _0966_ _1214_ _1216_ _0970_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3097_ _1146_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3999_ net47 _1414_ _1508_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Left_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_165_Left_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3020_ _0977_ _0999_ _1016_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_160_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_160_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4971_ clknet_leaf_38_clk _0303_ _0047_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3922_ _1882_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3853_ _0792_ _1823_ _0824_ _0781_ _0825_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_158_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2804_ _0851_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3784_ _1279_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2735_ net323 GCDdpath0.B_reg\[41\] VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2666_ _0715_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__or2_1
X_4405_ net346 _2262_ _2258_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__mux2_1
X_2597_ net312 GCDdpath0.B_reg\[31\] VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4336_ GCDdpath0.B_reg\[82\] net237 _2213_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4267_ _2165_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__clkbuf_1
X_3218_ _1136_ _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4198_ GCDdpath0.B_reg\[123\] net155 _2113_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__mux2_1
X_3149_ _1199_ GCDdpath0.B_reg\[36\] _0800_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2520_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5170_ clknet_leaf_5_clk _0502_ _0246_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dfrtp_4
X_4121_ net387 net128 _1406_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4052_ _0676_ _0677_ _1962_ _0680_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 operands_bits_A[102] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_3003_ _1048_ _1049_ _1050_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__or4b_1
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4954_ clknet_leaf_40_clk _0286_ _0030_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3905_ _1868_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4885_ _2456_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__inv_2
XFILLER_0_149_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3836_ _1807_ _1808_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3767_ _0709_ _1749_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2718_ _0762_ _0765_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__or3b_1
XFILLER_0_113_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3698_ _1326_ _1689_ _1690_ _1313_ GCDdpath0.B_reg\[69\] VGND VGND VPWR VPWR _1691_
+ sky130_fd_sc_hd__o32a_1
Xoutput330 net330 VGND VGND VPWR VPWR result_bits_data[48] sky130_fd_sc_hd__clkbuf_4
X_2649_ _0656_ _0659_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput341 net341 VGND VGND VPWR VPWR result_bits_data[58] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput352 net352 VGND VGND VPWR VPWR result_bits_data[68] sky130_fd_sc_hd__buf_2
Xoutput363 net363 VGND VGND VPWR VPWR result_bits_data[78] sky130_fd_sc_hd__clkbuf_4
Xoutput374 net374 VGND VGND VPWR VPWR result_bits_data[88] sky130_fd_sc_hd__clkbuf_4
Xoutput385 net385 VGND VGND VPWR VPWR result_bits_data[98] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_39_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4319_ _2202_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4670_ _2421_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3621_ _1511_ _1573_ _1623_ _1624_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_116_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3552_ _1336_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_133_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2503_ GCDdpath0.B_reg\[99\] _0553_ GCDdpath0.B_reg\[97\] GCDdpath0.B_reg\[96\] VGND
+ VGND VPWR VPWR _0554_ sky130_fd_sc_hd__or4_1
XFILLER_0_45_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3483_ _0553_ _1504_ _1442_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5153_ clknet_leaf_10_clk _0485_ _0229_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4104_ net32 _2039_ _2029_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__mux2_1
X_5084_ clknet_leaf_36_clk _0416_ _0160_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4035_ _1511_ _1979_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4937_ clknet_leaf_48_clk _0269_ _0013_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4868_ _2453_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3819_ _0742_ _0743_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4799_ _2442_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ _1031_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4722_ _2426_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_170_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4653_ _2418_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 operands_bits_A[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
X_3604_ _1006_ _1573_ _1004_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 operands_bits_A[2] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_4584_ net387 _2388_ _2386_ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__mux2_1
Xinput62 operands_bits_A[3] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput73 operands_bits_A[4] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 operands_bits_A[5] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
XFILLER_0_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput95 operands_bits_A[6] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3535_ _0876_ _0873_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3466_ _1490_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_168_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3397_ GCDdpath0.B_reg\[110\] _1417_ _1418_ _1430_ _1387_ VGND VGND VPWR VPWR _1431_
+ sky130_fd_sc_hd__o221a_1
X_5136_ clknet_leaf_24_clk _0468_ _0212_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5067_ clknet_leaf_46_clk _0399_ _0143_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4018_ _0668_ _1964_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3320_ _1105_ _1106_ _1108_ _1361_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_106_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3251_ _1154_ _1297_ _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3182_ _0887_ _0890_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2966_ net268 GCDdpath0.B_reg\[107\] VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__and2b_1
XFILLER_0_174_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4705_ _2427_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2897_ net350 GCDdpath0.B_reg\[66\] VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__and2b_1
XFILLER_0_161_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4636_ _2413_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4567_ net293 _2376_ _2372_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3518_ _1386_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_90_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4498_ _2313_ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_34_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3449_ _1059_ _1475_ _1058_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_51_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5119_ clknet_leaf_22_clk _0451_ _0195_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_722 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput230 operands_bits_B[76] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_1
Xinput241 operands_bits_B[86] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_145_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput252 operands_bits_B[96] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_69_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2820_ GCDdpath0.B_reg\[89\] net375 VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2751_ GCDdpath0.B_reg\[36\] net317 VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2682_ net331 GCDdpath0.B_reg\[49\] VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4421_ _2274_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4352_ GCDdpath0.B_reg\[77\] net231 _2213_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_165_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ net284 _1293_ _1347_ _1308_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_165_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4283_ net385 _2176_ _2172_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__mux2_1
X_3234_ _1284_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _0980_ _1215_ _0971_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3096_ GCDdpath0.B_reg\[124\] net287 VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__and2b_1
XFILLER_0_167_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3998_ GCDdpath0.B_reg\[26\] _1409_ _1947_ _1412_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2949_ net382 GCDdpath0.B_reg\[95\] VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4619_ net257 VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4970_ clknet_leaf_37_clk _0302_ _0046_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3921_ _1878_ _1881_ _1340_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3852_ _0805_ _1822_ _0835_ _0834_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2803_ _0852_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3783_ _1509_ _1759_ _1762_ _1763_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2734_ _0783_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2665_ GCDdpath0.B_reg\[57\] net340 VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4404_ GCDdpath0.B_reg\[62\] net215 _2256_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__mux2_1
X_2596_ GCDdpath0.B_reg\[31\] net312 VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4335_ _2141_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__buf_2
X_4266_ net264 _2164_ _2158_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3217_ _1135_ _1137_ _1132_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4197_ _2116_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_1
X_3148_ net317 VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3079_ _1128_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4120_ _2053_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__clkbuf_1
X_4051_ _1993_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 operands_bits_A[103] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3002_ _1051_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4953_ clknet_leaf_38_clk _0285_ _0029_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3904_ net322 _1867_ _1841_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4884_ _2456_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3835_ _0733_ _0736_ _1806_ _0735_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3766_ net392 _0840_ _1748_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_144_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2717_ _0766_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nor2_1
X_3697_ _0969_ _0972_ _1676_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__and3b_1
XFILLER_0_113_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2648_ _0697_ _0698_ _0647_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a21oi_1
Xoutput320 net320 VGND VGND VPWR VPWR result_bits_data[39] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR result_bits_data[49] sky130_fd_sc_hd__buf_2
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput342 net342 VGND VGND VPWR VPWR result_bits_data[59] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput353 net353 VGND VGND VPWR VPWR result_bits_data[69] sky130_fd_sc_hd__buf_2
Xoutput364 net364 VGND VGND VPWR VPWR result_bits_data[79] sky130_fd_sc_hd__clkbuf_4
Xoutput375 net375 VGND VGND VPWR VPWR result_bits_data[89] sky130_fd_sc_hd__clkbuf_4
X_2579_ GCDdpath0.B_reg\[10\] net271 VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or2b_1
Xoutput386 net386 VGND VGND VPWR VPWR result_bits_data[99] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_39_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4318_ net374 _2200_ _2201_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4249_ net269 _2152_ _2144_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3620_ _0895_ _1313_ _1386_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3551_ GCDdpath0.B_reg\[89\] _1563_ _1482_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2502_ GCDdpath0.B_reg\[98\] VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3482_ _1047_ _1499_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5152_ clknet_leaf_12_clk _0484_ _0228_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4103_ GCDdpath0.B_reg\[12\] _2038_ _1989_ VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__mux2_1
X_5083_ clknet_leaf_35_clk _0415_ _0159_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4034_ _0671_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4936_ clknet_leaf_47_clk _0268_ _0012_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_10 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4867_ _2453_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3818_ _1322_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__buf_2
XFILLER_0_160_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4798_ _2442_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3749_ net87 _1506_ _1734_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2982_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4721_ _2429_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4652_ _2418_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput30 operands_bits_A[126] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3603_ _0571_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput41 operands_bits_A[20] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput52 operands_bits_A[30] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
X_4583_ GCDdpath0.B_reg\[9\] net256 _2384_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__mux2_1
Xinput63 operands_bits_A[40] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
Xinput74 operands_bits_A[50] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 operands_bits_A[60] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
X_3534_ _1326_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput96 operands_bits_A[70] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_149_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3465_ net262 _1488_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3396_ _1034_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__xnor2_1
X_5135_ clknet_leaf_14_clk _0467_ _0211_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5066_ clknet_leaf_43_clk _0398_ _0142_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4017_ _0686_ _0688_ _1963_ _0687_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__o31a_1
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4919_ _2461_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3250_ _1299_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3181_ _1229_ _1231_ _0886_ _0882_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2965_ _1000_ _0853_ _1002_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4704_ _2427_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2896_ GCDdpath0.B_reg\[66\] net350 VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4635_ _2415_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ GCDdpath0.B_reg\[14\] net162 _2370_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3517_ _0854_ _1530_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4497_ _2327_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3448_ _1066_ _1474_ _1065_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _1302_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__buf_2
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5118_ clknet_leaf_24_clk _0450_ _0194_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5049_ clknet_leaf_49_clk _0381_ _0125_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput220 operands_bits_B[67] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput231 operands_bits_B[77] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput242 operands_bits_B[87] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_145_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput253 operands_bits_B[97] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_106_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2750_ _0799_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2681_ net330 GCDdpath0.B_reg\[48\] VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4420_ net392 _2271_ _2273_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4351_ _2224_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3302_ GCDdpath0.B_reg\[121\] _1313_ _1343_ _1346_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _0553_ net254 _2170_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _1277_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3164_ _0952_ _0955_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3095_ net287 GCDdpath0.B_reg\[124\] VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3997_ _1343_ _1940_ _1946_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__nor3_1
XFILLER_0_174_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2948_ _0912_ _0998_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2879_ _0926_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4618_ _2409_ _1408_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4549_ GCDdpath0.B_reg\[19\] net167 _2356_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3920_ GCDdpath0.B_reg\[37\] _1880_ _1834_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3851_ _0769_ _1821_ _0818_ _0822_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2802_ GCDdpath0.B_reg\[94\] net381 VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__or2b_1
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3782_ GCDdpath0.B_reg\[57\] _1516_ _1517_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2733_ GCDdpath0.B_reg\[42\] net324 VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2664_ net340 GCDdpath0.B_reg\[57\] VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4403_ _2261_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
X_2595_ _0642_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_97_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4334_ _2212_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4265_ GCDdpath0.B_reg\[103\] net133 _2156_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__mux2_1
X_3216_ _1128_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__inv_2
X_4196_ net287 _2114_ _2115_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3147_ _0821_ _1196_ _1197_ _0805_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a31o_1
X_3078_ GCDdpath0.B_reg\[123\] net286 VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4050_ net298 _1991_ _1992_ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3001_ GCDdpath0.B_reg\[96\] net383 VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__and2b_1
Xinput6 operands_bits_A[104] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4952_ clknet_leaf_40_clk _0284_ _0028_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3903_ net63 _1866_ _1817_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4883_ _2456_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3834_ _0733_ _0735_ _0736_ _1806_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_138_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3765_ _0839_ _1747_ _0710_ _0715_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2716_ net314 GCDdpath0.B_reg\[33\] VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3696_ _0972_ _1676_ _0969_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput310 net310 VGND VGND VPWR VPWR result_bits_data[2] sky130_fd_sc_hd__clkbuf_4
X_2647_ GCDdpath0.B_reg\[30\] net311 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__and2b_1
Xoutput321 net321 VGND VGND VPWR VPWR result_bits_data[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput332 net332 VGND VGND VPWR VPWR result_bits_data[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput343 net343 VGND VGND VPWR VPWR result_bits_data[5] sky130_fd_sc_hd__clkbuf_4
Xoutput354 net354 VGND VGND VPWR VPWR result_bits_data[6] sky130_fd_sc_hd__clkbuf_4
X_2578_ net282 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__inv_2
Xoutput365 net365 VGND VGND VPWR VPWR result_bits_data[7] sky130_fd_sc_hd__clkbuf_4
Xoutput376 net376 VGND VGND VPWR VPWR result_bits_data[8] sky130_fd_sc_hd__clkbuf_4
Xoutput387 net387 VGND VGND VPWR VPWR result_bits_data[9] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_39_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4317_ _2186_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__buf_2
X_4248_ GCDdpath0.B_reg\[108\] net138 _2142_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__mux2_1
X_4179_ net394 GCDdpath0.B_reg\[0\] VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3550_ _1561_ _1562_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2501_ GCDdpath0.B_reg\[111\] GCDdpath0.B_reg\[110\] GCDdpath0.B_reg\[109\] GCDdpath0.B_reg\[108\]
+ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or4_1
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3481_ _1354_ _1497_ _1503_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5151_ clknet_leaf_9_clk _0483_ _0227_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4102_ _2018_ _2037_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5082_ clknet_leaf_39_clk _0414_ _0158_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4033_ _0693_ _0536_ _1965_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4935_ clknet_leaf_47_clk _0267_ _0011_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 net357 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4866_ _2453_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3817_ net335 _1294_ _1792_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__o21a_1
X_4797_ _2442_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3748_ _0515_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3679_ _0956_ _1673_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__or2_2
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2981_ net272 GCDdpath0.B_reg\[110\] VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4720_ _2429_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_170_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4651_ _2418_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 operands_bits_A[117] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ net110 _1341_ _1342_ _1608_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__o31a_1
Xinput31 operands_bits_A[127] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
X_4582_ _2387_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 operands_bits_A[21] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput53 operands_bits_A[31] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput64 operands_bits_A[41] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xinput75 operands_bits_A[51] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
X_3533_ _1548_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_1
Xinput86 operands_bits_A[61] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 operands_bits_A[71] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3464_ _1292_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3395_ _1082_ _1424_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5134_ clknet_leaf_15_clk _0466_ _0210_ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dfrtp_4
X_5065_ clknet_leaf_46_clk _0397_ _0141_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4016_ _0676_ _0677_ _1962_ _0680_ _0673_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_168_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4918_ _2461_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_33_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4849_ _2450_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3180_ _1003_ _1230_ _0883_ _0900_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__a211o_1
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2964_ _0879_ _1012_ _1014_ _0862_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__o22a_1
XFILLER_0_158_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4703_ _2427_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2895_ _0944_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4634_ _2415_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4565_ _2375_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3516_ net382 _1445_ _1533_ _1534_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4496_ net316 _2326_ _2316_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ _1063_ _1473_ _1062_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _1406_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__buf_2
X_5117_ clknet_leaf_24_clk _0449_ _0193_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5048_ clknet_leaf_1_clk _0380_ _0124_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_108_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput210 operands_bits_B[58] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
Xinput221 operands_bits_B[68] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
Xinput232 operands_bits_B[78] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput243 operands_bits_B[88] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput254 operands_bits_B[98] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_106_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2680_ _0718_ _0724_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4350_ net363 _2223_ _2215_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3301_ _1344_ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__xnor2_1
X_4281_ _2175_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_165_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3232_ _1158_ _0575_ _1154_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_3_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_3163_ _0944_ _0978_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3094_ net288 GCDdpath0.B_reg\[125\] VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3996_ _0641_ _1939_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ _0942_ _0986_ _0992_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_44_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2878_ _0927_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4617_ _2409_ _2411_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4548_ _2363_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4479_ GCDdpath0.B_reg\[40\] net191 _2314_ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_160_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3850_ _0684_ _0708_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2801_ net381 GCDdpath0.B_reg\[94\] VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__or2b_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3781_ _1511_ _1761_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2732_ net324 GCDdpath0.B_reg\[42\] VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2663_ _0712_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4402_ net347 _2260_ _2258_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2594_ _0643_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4333_ net369 _2211_ _2201_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__mux2_1
X_4264_ _2163_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3215_ _1124_ _1265_ _1100_ _1105_ _1107_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__a2111oi_1
XPHY_EDGE_ROW_163_Right_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4195_ _2082_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__buf_2
XFILLER_0_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3146_ net315 _0819_ GCDdpath0.B_reg\[34\] VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3077_ net286 GCDdpath0.B_reg\[123\] VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3979_ _1928_ _1931_ _1340_ VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3000_ net383 GCDdpath0.B_reg\[96\] VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 operands_bits_A[105] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4951_ clknet_leaf_41_clk _0283_ _0027_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3902_ GCDdpath0.B_reg\[40\] _1865_ _1810_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4882_ _2456_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3833_ _0837_ _1722_ _1770_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_138_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3764_ _0714_ _1724_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2715_ GCDdpath0.B_reg\[33\] net314 VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3695_ _1688_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput300 net300 VGND VGND VPWR VPWR result_bits_data[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2646_ _0648_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__inv_2
Xoutput311 net311 VGND VGND VPWR VPWR result_bits_data[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput322 net322 VGND VGND VPWR VPWR result_bits_data[40] sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR result_bits_data[50] sky130_fd_sc_hd__buf_2
XFILLER_0_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput344 net344 VGND VGND VPWR VPWR result_bits_data[60] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2577_ _0609_ _0611_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput355 net355 VGND VGND VPWR VPWR result_bits_data[70] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput366 net366 VGND VGND VPWR VPWR result_bits_data[80] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput377 net377 VGND VGND VPWR VPWR result_bits_data[90] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput388 net388 VGND VGND VPWR VPWR result_val sky130_fd_sc_hd__clkbuf_4
X_4316_ GCDdpath0.B_reg\[88\] net243 _2199_ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4247_ _2151_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__clkbuf_1
X_4178_ net299 _1407_ _2101_ _2102_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3129_ _0743_ _0740_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__or2b_1
XFILLER_0_167_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2500_ GCDdpath0.B_reg\[107\] GCDdpath0.B_reg\[106\] GCDdpath0.B_reg\[105\] GCDdpath0.B_reg\[104\]
+ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3480_ GCDdpath0.B_reg\[99\] _1325_ _1409_ _1502_ _1415_ VGND VGND VPWR VPWR _1503_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5150_ clknet_leaf_12_clk _0482_ _0226_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4101_ _0617_ _2017_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__nor2_1
X_5081_ clknet_leaf_38_clk _0413_ _0157_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dfrtp_4
X_4032_ net301 net42 _1406_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4934_ clknet_leaf_48_clk _0266_ _0010_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4865_ _2447_ VGND VGND VPWR VPWR _2453_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 net361 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_170_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3816_ net76 _1609_ _1790_ _1791_ _1407_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4796_ _2442_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3747_ GCDdpath0.B_reg\[62\] _1732_ _1442_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3678_ _0808_ _0848_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2629_ net296 GCDdpath0.B_reg\[17\] VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_93_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ GCDdpath0.B_reg\[110\] net272 VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_174_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4650_ _2413_ VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 operands_bits_A[108] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_3601_ net369 _1539_ _1607_ _1306_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__o22a_1
XFILLER_0_142_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput21 operands_bits_A[118] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput32 operands_bits_A[12] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
X_4581_ net271 _2385_ _2386_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__mux2_1
Xinput43 operands_bits_A[22] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput54 operands_bits_A[32] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput65 operands_bits_A[42] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
X_3532_ net379 _1547_ _1489_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__mux2_1
Xinput76 operands_bits_A[52] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput87 operands_bits_A[62] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
Xinput98 operands_bits_A[72] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3463_ net3 _1487_ _1468_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3394_ net273 _1324_ _1427_ _1428_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5133_ clknet_leaf_18_clk _0465_ _0209_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dfrtp_4
X_5064_ clknet_leaf_0_clk _0396_ _0140_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4015_ _1961_ _1174_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__nand2_2
XFILLER_0_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4917_ _2461_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4848_ _2450_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4779_ _2433_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_160_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2963_ _0866_ GCDdpath0.B_reg\[90\] _0863_ _0864_ _1013_ VGND VGND VPWR VPWR _1014_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4702_ _2427_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2894_ _0943_ _0564_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4633_ _2415_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4564_ net294 _2374_ _2372_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3515_ net123 _1432_ _1479_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__o21a_1
X_4495_ GCDdpath0.B_reg\[35\] net185 _2314_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3446_ _1472_ _1421_ _1076_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_51_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ GCDdpath0.B_reg\[112\] _1409_ _1411_ _1412_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__a211o_1
X_5116_ clknet_leaf_23_clk _0448_ _0192_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dfrtp_4
X_5047_ clknet_leaf_1_clk _0379_ _0123_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput200 operands_bits_B[49] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_1
Xinput211 operands_bits_B[59] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
Xinput222 operands_bits_B[69] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
Xinput233 operands_bits_B[79] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput244 operands_bits_B[89] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput255 operands_bits_B[99] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_106_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3300_ _1138_ _1328_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__and2b_1
X_4280_ net386 _2174_ _2172_ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_165_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _1281_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__buf_2
X_3162_ _1179_ _1185_ _1211_ _1212_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_55_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3093_ _1134_ _1135_ _1142_ _1143_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3995_ net307 _1293_ _1944_ _0573_ _1945_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2946_ _0993_ _0935_ _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2877_ net361 GCDdpath0.B_reg\[76\] VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4616_ _0518_ _0543_ _0568_ net258 _2410_ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__o32a_1
XFILLER_0_103_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4547_ net300 _2362_ _2358_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4478_ _2313_ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3429_ _1023_ _1024_ _1447_ _1025_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_5_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2800_ _0849_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_158_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3780_ _0717_ _1760_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2731_ _0780_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2662_ GCDdpath0.B_reg\[56\] net339 VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_136_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4401_ GCDdpath0.B_reg\[63\] net216 _2256_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2593_ net305 GCDdpath0.B_reg\[25\] VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4332_ GCDdpath0.B_reg\[83\] net238 _2199_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4263_ net265 _2162_ _2158_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3214_ _1094_ _1101_ _1263_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__or4_1
X_4194_ GCDdpath0.B_reg\[124\] net156 _2113_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3145_ _0764_ _1195_ _0766_ _0762_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3076_ _1105_ _1119_ _1126_ _1110_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__o22a_1
XFILLER_0_167_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3978_ GCDdpath0.B_reg\[29\] _1930_ _1834_ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__mux2_1
X_2929_ _0943_ _0564_ _0948_ _0951_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 operands_bits_A[106] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4950_ clknet_leaf_41_clk _0282_ _0026_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3901_ _1863_ _1864_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4881_ _2456_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3832_ net333 _1793_ _1803_ _1559_ _1805_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3763_ _1746_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2714_ _0763_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or2b_1
XFILLER_0_125_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3694_ net355 _1686_ _1687_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2645_ _0690_ _0692_ _0695_ _0663_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a31o_1
Xoutput301 net301 VGND VGND VPWR VPWR result_bits_data[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput312 net312 VGND VGND VPWR VPWR result_bits_data[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput323 net323 VGND VGND VPWR VPWR result_bits_data[41] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput334 net334 VGND VGND VPWR VPWR result_bits_data[51] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2576_ net292 _0625_ _0615_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a21o_1
Xoutput345 net345 VGND VGND VPWR VPWR result_bits_data[61] sky130_fd_sc_hd__buf_2
XFILLER_0_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput356 net356 VGND VGND VPWR VPWR result_bits_data[71] sky130_fd_sc_hd__buf_2
Xoutput367 net367 VGND VGND VPWR VPWR result_bits_data[81] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput378 net378 VGND VGND VPWR VPWR result_bits_data[91] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4315_ _2141_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4246_ net270 _2150_ _2144_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__mux2_1
X_4177_ net40 _1496_ _1508_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3128_ _1167_ _1173_ _1178_ _0807_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__a31oi_2
XPHY_EDGE_ROW_153_Left_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3059_ _1105_ _1106_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__or3_1
XFILLER_0_167_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Left_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_171_Left_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4100_ _2036_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5080_ clknet_leaf_40_clk _0412_ _0156_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dfrtp_4
X_4031_ net393 _1408_ _1975_ _1976_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4933_ clknet_leaf_48_clk _0265_ _0009_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4864_ _2452_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_13 net363 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3815_ GCDdpath0.B_reg\[52\] _1281_ _1386_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4795_ _2442_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3746_ _0722_ _1727_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3677_ _1672_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2628_ net295 GCDdpath0.B_reg\[16\] VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2559_ _0608_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4229_ _2138_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3600_ _1300_ _1605_ _1606_ _1313_ GCDdpath0.B_reg\[83\] VGND VGND VPWR VPWR _1607_
+ sky130_fd_sc_hd__o32a_1
Xinput11 operands_bits_A[109] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 operands_bits_A[119] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
X_4580_ _1295_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput33 operands_bits_A[13] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput44 operands_bits_A[23] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput55 operands_bits_A[33] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
X_3531_ net120 _1546_ _1468_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__mux2_1
Xinput66 operands_bits_A[43] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput77 operands_bits_A[53] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
XFILLER_0_80_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput88 operands_bits_A[63] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput99 operands_bits_A[73] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_1
X_3462_ GCDdpath0.B_reg\[101\] _1486_ _1482_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3393_ net14 _1305_ _1369_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5132_ clknet_leaf_18_clk _0464_ _0208_ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dfrtp_4
X_5063_ clknet_leaf_47_clk _0395_ _0139_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4014_ _1960_ _0679_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4916_ _2461_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4847_ _2450_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4778_ _2438_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3729_ _1280_ _1674_ _1715_ _1716_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_724 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2962_ _0870_ _0875_ _0874_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__or3b_1
XFILLER_0_158_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4701_ _2426_ VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2893_ _0943_ _0564_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__nand2_2
XFILLER_0_173_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4632_ _2415_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4563_ GCDdpath0.B_reg\[15\] net163 _2370_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3514_ GCDdpath0.B_reg\[95\] _1417_ _1418_ _1532_ _1387_ VGND VGND VPWR VPWR _1533_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_142_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4494_ _2325_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3445_ _1054_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _0571_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ clknet_leaf_23_clk _0447_ _0191_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5046_ clknet_leaf_49_clk _0378_ _0122_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput201 operands_bits_B[4] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
Xinput212 operands_bits_B[5] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput223 operands_bits_B[6] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
Xinput234 operands_bits_B[7] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 operands_bits_B[8] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_145_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput256 operands_bits_B[9] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_106_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3230_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__buf_2
X_3161_ _1070_ _0912_ _0976_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__nor3_2
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3092_ _1128_ _1132_ _1129_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3994_ net48 _1804_ _0516_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2945_ _0993_ _0937_ _0995_ _0932_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2876_ GCDdpath0.B_reg\[76\] net361 VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4615_ net388 VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4546_ _0536_ net169 _2356_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4477_ _1404_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__buf_2
X_3428_ _1457_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__clkbuf_1
X_3359_ _1071_ _1092_ _1115_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_5_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ clknet_leaf_8_clk _0361_ _0105_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2730_ GCDdpath0.B_reg\[43\] net325 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2661_ net339 GCDdpath0.B_reg\[56\] VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_136_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4400_ _2259_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2592_ GCDdpath0.B_reg\[25\] net305 VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4331_ _2210_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4262_ GCDdpath0.B_reg\[104\] net134 _2156_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3213_ _1093_ _1095_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4193_ _1405_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_66_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3144_ net314 GCDdpath0.B_reg\[33\] VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__or2b_1
XFILLER_0_158_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3075_ _1104_ _1123_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__o21a_1
XFILLER_0_173_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_166_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3977_ _0661_ _1929_ VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_75_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2928_ _0944_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _0898_ _0901_ _0904_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4529_ GCDdpath0.B_reg\[25\] net174 _2342_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput9 operands_bits_A[107] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3900_ _0791_ _1823_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4880_ _2454_ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3831_ net74 _1804_ _1734_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_138_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3762_ net344 _1744_ _1745_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2713_ net313 GCDdpath0.B_reg\[32\] VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__or2b_1
X_3693_ _1601_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2644_ _0664_ _0667_ _0669_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput302 net393 VGND VGND VPWR VPWR result_bits_data[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput313 net313 VGND VGND VPWR VPWR result_bits_data[32] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput324 net324 VGND VGND VPWR VPWR result_bits_data[42] sky130_fd_sc_hd__buf_2
XFILLER_0_125_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2575_ net292 _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or2_1
Xoutput335 net335 VGND VGND VPWR VPWR result_bits_data[52] sky130_fd_sc_hd__buf_2
XFILLER_0_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput346 net346 VGND VGND VPWR VPWR result_bits_data[62] sky130_fd_sc_hd__buf_2
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput357 net357 VGND VGND VPWR VPWR result_bits_data[72] sky130_fd_sc_hd__buf_2
Xoutput368 net368 VGND VGND VPWR VPWR result_bits_data[82] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4314_ _2198_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput379 net379 VGND VGND VPWR VPWR result_bits_data[92] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4245_ GCDdpath0.B_reg\[109\] net139 _2142_ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__mux2_1
X_4176_ GCDdpath0.B_reg\[1\] _1327_ _2100_ _1412_ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__a211o_1
X_3127_ _0683_ _1174_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_171_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3058_ _1107_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4030_ net43 _1414_ _1508_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4932_ clknet_leaf_0_clk _0264_ _0008_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[5\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_44_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4863_ _2452_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_14 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3814_ _1773_ _1789_ _1296_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4794_ _2440_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3745_ net347 _1349_ _1730_ _1731_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o22a_1
XFILLER_0_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3676_ net357 _1671_ _1602_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2627_ _0676_ _0677_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2558_ GCDdpath0.B_reg\[9\] net387 VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2489_ GCDdpath0.B_reg\[19\] GCDdpath0.B_reg\[18\] GCDdpath0.B_reg\[17\] GCDdpath0.B_reg\[16\]
+ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_54_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4228_ net276 _2137_ _2129_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4159_ _1395_ _2066_ _2085_ _2086_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout392 net341 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_21_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput12 operands_bits_A[10] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput23 operands_bits_A[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput34 operands_bits_A[14] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
XFILLER_0_108_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput45 operands_bits_A[24] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3530_ GCDdpath0.B_reg\[92\] _1545_ _1482_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput56 operands_bits_A[34] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput67 operands_bits_A[44] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput78 operands_bits_A[54] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xinput89 operands_bits_A[64] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlymetal6s2s_1
X_3461_ _1067_ _1474_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3392_ GCDdpath0.B_reg\[111\] _1417_ _1418_ _1426_ _1387_ VGND VGND VPWR VPWR _1427_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5131_ clknet_leaf_18_clk _0463_ _0207_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dfrtp_4
X_5062_ clknet_leaf_48_clk _0394_ _0138_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4013_ GCDdpath0.B_reg\[16\] net295 VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4915_ _2408_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4846_ _2450_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ _2438_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3728_ GCDdpath0.B_reg\[64\] _1520_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3659_ _1222_ _1652_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2961_ _0894_ _1008_ _1009_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4700_ _2408_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__buf_2
XFILLER_0_173_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2892_ net351 VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4631_ _2415_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4562_ _2373_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3513_ _0851_ _1531_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__xnor2_1
X_4493_ net317 _2324_ _2316_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_3444_ _1056_ _1057_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3375_ _1343_ _1396_ _1410_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5114_ clknet_leaf_14_clk _0446_ _0190_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5045_ clknet_leaf_49_clk _0377_ _0121_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4829_ reset VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput202 operands_bits_B[50] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput213 operands_bits_B[60] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput224 operands_bits_B[70] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
Xinput235 operands_bits_B[80] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 operands_bits_B[90] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput257 operands_val VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
XFILLER_0_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3160_ _0719_ _1192_ _1210_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__o21ai_2
Xhold1 GCDdpath0.B_reg\[71\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _1136_ _1138_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3993_ GCDdpath0.B_reg\[27\] _1943_ _1281_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2944_ _0925_ _0927_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2875_ _0924_ _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4614_ _2408_ VGND VGND VPWR VPWR _2409_ sky130_fd_sc_hd__buf_2
XFILLER_0_115_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4545_ _2361_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4476_ _2312_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3427_ net267 _1456_ _1393_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3358_ _1279_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__clkbuf_4
X_3289_ GCDdpath0.B_reg\[122\] _1334_ _1319_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux2_1
X_5028_ clknet_leaf_9_clk _0360_ _0104_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2660_ _0709_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2591_ _0639_ _0640_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4330_ net370 _2209_ _2201_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4261_ _2161_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3212_ _1112_ _1114_ _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4192_ _2112_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3143_ _0782_ _0785_ _1193_ _0787_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_2_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3074_ _1100_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_783 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ _0656_ _1917_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2927_ _0943_ GCDdpath0.B_reg\[67\] _0947_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2858_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2789_ GCDdpath0.B_reg\[58\] VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4528_ _2349_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4459_ _2272_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3830_ _1302_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__buf_2
XFILLER_0_157_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3761_ _1601_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2712_ GCDdpath0.B_reg\[32\] net313 VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3692_ net96 _1685_ _1665_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2643_ _0693_ _0536_ _0670_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput303 net303 VGND VGND VPWR VPWR result_bits_data[23] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput314 net314 VGND VGND VPWR VPWR result_bits_data[33] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput325 net325 VGND VGND VPWR VPWR result_bits_data[43] sky130_fd_sc_hd__clkbuf_4
X_2574_ GCDdpath0.B_reg\[13\] VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__inv_2
Xoutput336 net336 VGND VGND VPWR VPWR result_bits_data[53] sky130_fd_sc_hd__buf_2
XFILLER_0_65_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput347 net347 VGND VGND VPWR VPWR result_bits_data[63] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput358 net358 VGND VGND VPWR VPWR result_bits_data[73] sky130_fd_sc_hd__buf_2
X_4313_ net375 _2197_ _2187_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput369 net369 VGND VGND VPWR VPWR result_bits_data[83] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4244_ _2149_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_1
X_4175_ _0582_ _1620_ _2099_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__and3_1
X_3126_ _0683_ _0623_ _0598_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__nor4_1
XFILLER_0_171_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3057_ GCDdpath0.B_reg\[118\] net280 VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3959_ _0624_ _0638_ _0682_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4931_ clknet_leaf_0_clk _0263_ _0007_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4862_ _2452_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3813_ _0756_ _1788_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_15 net388 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_172_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4793_ _2441_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3744_ net88 _1583_ _1517_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3675_ net98 _1670_ _1665_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2626_ GCDdpath0.B_reg\[17\] net296 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_101_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2557_ net387 GCDdpath0.B_reg\[9\] VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2488_ GCDdpath0.B_reg\[31\] GCDdpath0.B_reg\[30\] GCDdpath0.B_reg\[29\] GCDdpath0.B_reg\[28\]
+ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or4_1
X_4227_ GCDdpath0.B_reg\[114\] net145 _2127_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4158_ GCDdpath0.B_reg\[4\] _1398_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__and2_1
X_3109_ net297 _0688_ GCDdpath0.B_reg\[18\] VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__or3b_1
X_4089_ GCDdpath0.B_reg\[14\] _1299_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout393 net302 VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 operands_bits_A[110] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput24 operands_bits_A[120] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 operands_bits_A[15] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
XFILLER_0_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput46 operands_bits_A[25] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 operands_bits_A[35] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
Xinput68 operands_bits_A[45] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput79 operands_bits_A[55] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_172_Right_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3460_ _1485_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3391_ _1419_ _1425_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5130_ clknet_leaf_20_clk _0462_ _0206_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_36_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5061_ clknet_leaf_48_clk _0393_ _0137_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dfrtp_4
X_4012_ _1959_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4914_ _2460_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4845_ _2450_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4776_ _2438_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3727_ _0956_ _1673_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3658_ net360 _1440_ _1655_ _1559_ _1656_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2609_ net309 GCDdpath0.B_reg\[29\] VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3589_ _1577_ _1596_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Left_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_168_Left_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2960_ net372 _1010_ _0891_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_174_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2891_ _0923_ _0931_ _0938_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__or4_1
XFILLER_0_139_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4630_ _2415_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4561_ net295 _2371_ _2372_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3512_ _0852_ _1530_ _0853_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__a21bo_1
X_4492_ GCDdpath0.B_reg\[36\] net186 _2314_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3443_ _1470_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3374_ _1115_ _1071_ _1092_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5113_ clknet_leaf_14_clk _0445_ _0189_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_51_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5044_ clknet_leaf_49_clk _0376_ _0120_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4828_ _2446_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4759_ _2436_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput203 operands_bits_B[51] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
Xinput214 operands_bits_B[61] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput225 operands_bits_B[71] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput236 operands_bits_B[81] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 operands_bits_B[91] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_145_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 result_rdy VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_162_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 net260 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _1118_ _1127_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3992_ _1941_ _1942_ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2943_ GCDdpath0.B_reg\[77\] net362 VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__and2b_1
XFILLER_0_174_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2874_ net362 GCDdpath0.B_reg\[77\] VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__or2b_2
XTAP_TAPCELL_ROW_44_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4613_ reset VGND VGND VPWR VPWR _2408_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4544_ net301 _2360_ _2358_ VGND VGND VPWR VPWR _2361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4475_ net323 _2311_ _2301_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3426_ net8 _1455_ _1337_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3357_ _1394_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__clkbuf_1
X_3288_ _1133_ _1329_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__xnor2_1
X_5027_ clknet_leaf_9_clk _0359_ _0103_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_68_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2590_ net306 GCDdpath0.B_reg\[26\] VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4260_ net266 _2160_ _2158_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3211_ _1098_ _1111_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nor2_1
X_4191_ net288 _2111_ _1282_ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3142_ _0786_ _0789_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3073_ _1099_ _1102_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3975_ net309 net50 _1615_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2926_ _0808_ _0848_ _0912_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2857_ _0906_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2788_ _0713_ _0716_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4527_ net306 _2348_ _2344_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4458_ _0526_ net197 _2299_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__mux2_1
X_3409_ _1041_ _1423_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__xor2_1
X_4389_ _2251_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_123_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3760_ net85 _1743_ _1718_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2711_ _0760_ _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3691_ GCDdpath0.B_reg\[70\] _1683_ _1684_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2642_ net300 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput304 net304 VGND VGND VPWR VPWR result_bits_data[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput315 net315 VGND VGND VPWR VPWR result_bits_data[34] sky130_fd_sc_hd__clkbuf_4
X_2573_ _0599_ _0601_ _0604_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a31o_1
Xoutput326 net326 VGND VGND VPWR VPWR result_bits_data[44] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput337 net337 VGND VGND VPWR VPWR result_bits_data[54] sky130_fd_sc_hd__clkbuf_4
X_4312_ GCDdpath0.B_reg\[89\] net244 _2184_ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput348 net348 VGND VGND VPWR VPWR result_bits_data[64] sky130_fd_sc_hd__clkbuf_4
Xoutput359 net359 VGND VGND VPWR VPWR result_bits_data[74] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4243_ net272 _2148_ _2144_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4174_ net394 _0580_ _0581_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__or3_1
X_3125_ net394 _0580_ _0584_ _0582_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_171_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3056_ net280 GCDdpath0.B_reg\[118\] VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3958_ _0647_ _0648_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2909_ _0958_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3889_ GCDdpath0.B_reg\[42\] _1854_ _1810_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_131_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_140_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4930_ clknet_leaf_0_clk _0262_ _0006_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4861_ _2452_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3812_ _0810_ _1772_ _0742_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__a21o_1
X_4792_ _2441_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
XANTENNA_16 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3743_ GCDdpath0.B_reg\[63\] _1285_ _1549_ _1729_ _1536_ VGND VGND VPWR VPWR _1730_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3674_ GCDdpath0.B_reg\[72\] _1669_ _1598_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2625_ GCDdpath0.B_reg\[16\] net295 VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2556_ _0605_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2487_ GCDdpath0.B_reg\[27\] GCDdpath0.B_reg\[26\] GCDdpath0.B_reg\[25\] GCDdpath0.B_reg\[24\]
+ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4226_ _2136_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4157_ _0597_ _2065_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__nand2_1
X_3108_ _0576_ _1154_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a21bo_1
X_4088_ _0605_ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3039_ _1082_ _1041_ _1087_ _1088_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__o311a_1
XFILLER_0_167_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout394 net260 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 operands_bits_A[111] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput25 operands_bits_A[121] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
XFILLER_0_154_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput36 operands_bits_A[16] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput47 operands_bits_A[26] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xinput58 operands_bits_A[36] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 operands_bits_A[46] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3390_ _1032_ _1082_ _1424_ _1031_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__o31a_1
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5060_ clknet_leaf_0_clk _0392_ _0136_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dfrtp_4
X_4011_ net304 _1958_ _1911_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4913_ _2460_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4844_ _2447_ VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4775_ _2438_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3726_ net349 _1408_ _1713_ _1714_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3657_ net101 _1506_ _1355_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2608_ GCDdpath0.B_reg\[29\] net309 VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_73_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3588_ _1575_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2539_ net354 GCDdpath0.B_reg\[6\] VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4209_ _2124_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2890_ _0939_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4560_ _1295_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3511_ _1525_ _1529_ _0859_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__o21ba_1
X_4491_ _2323_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
X_3442_ net265 _1469_ _1393_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3373_ _1300_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ clknet_leaf_39_clk _0444_ _0188_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_51_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5043_ clknet_leaf_48_clk _0375_ _0119_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4827_ _2446_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4758_ _2433_ VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3709_ _0947_ _1675_ _0946_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__o21ai_1
X_4689_ _2424_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput204 operands_bits_B[52] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
Xinput215 operands_bits_B[62] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
Xinput226 operands_bits_B[72] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_1
Xinput237 operands_bits_B[82] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_145_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 operands_bits_B[92] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_145_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3 net259 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3991_ _0639_ _0640_ _0703_ _1940_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2942_ _0933_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2873_ GCDdpath0.B_reg\[77\] net362 VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_44_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4612_ _2407_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4543_ GCDdpath0.B_reg\[21\] net170 _2356_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4474_ GCDdpath0.B_reg\[41\] net192 _2299_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__mux2_1
X_3425_ GCDdpath0.B_reg\[106\] _1454_ _1319_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3356_ net276 _1392_ _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3287_ net286 _1324_ _1332_ _1333_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5026_ clknet_leaf_10_clk _0358_ _0102_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_68_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3210_ _1105_ _1108_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__and2b_1
X_4190_ GCDdpath0.B_reg\[125\] net157 _1904_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3141_ _0720_ _1186_ _1191_ _0721_ _0723_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__o311a_1
XFILLER_0_158_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_174_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3072_ _1098_ _1120_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_167_Right_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3974_ net311 _1793_ _1926_ _0573_ _1927_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_63_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2925_ _0942_ _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__or2b_2
XFILLER_0_45_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2856_ _0905_ GCDdpath0.B_reg\[82\] VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2787_ _0727_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__inv_2
X_4526_ GCDdpath0.B_reg\[26\] net175 _2342_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4457_ _2227_ VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__buf_2
XFILLER_0_141_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3408_ _1322_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4388_ net351 _2250_ _2244_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__mux2_1
X_3339_ GCDdpath0.B_reg\[116\] _1378_ _1319_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5009_ clknet_leaf_15_clk _0341_ _0085_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2710_ net315 GCDdpath0.B_reg\[34\] VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__xor2_2
XFILLER_0_171_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3690_ _1318_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__buf_2
X_2641_ net393 _0691_ _0666_ _0665_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput305 net305 VGND VGND VPWR VPWR result_bits_data[25] sky130_fd_sc_hd__clkbuf_4
X_2572_ _0607_ _0614_ _0619_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or4_1
XFILLER_0_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput316 net316 VGND VGND VPWR VPWR result_bits_data[35] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput327 net327 VGND VGND VPWR VPWR result_bits_data[45] sky130_fd_sc_hd__buf_2
Xoutput338 net338 VGND VGND VPWR VPWR result_bits_data[55] sky130_fd_sc_hd__buf_2
X_4311_ _2196_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__clkbuf_1
Xoutput349 net349 VGND VGND VPWR VPWR result_bits_data[65] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4242_ GCDdpath0.B_reg\[110\] net141 _2142_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__mux2_1
X_4173_ net310 _1407_ _2097_ _2098_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__a22o_1
X_3124_ _0587_ _0586_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3055_ GCDdpath0.B_reg\[119\] net281 VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_47_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3957_ _1912_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2908_ GCDdpath0.B_reg\[70\] net355 VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3888_ _0785_ _1853_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2839_ net373 GCDdpath0.B_reg\[87\] VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4509_ GCDdpath0.B_reg\[31\] net181 _2328_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_38_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_159_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_172_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4860_ _2452_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3811_ net77 _1415_ _0517_ _1787_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o31a_1
XFILLER_0_172_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4791_ _2441_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 net353 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3742_ _1721_ _1728_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__xor2_1
XFILLER_0_172_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3673_ _1628_ _1668_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2624_ _0673_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2555_ net294 GCDdpath0.B_reg\[15\] VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_93_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2486_ GCDdpath0.B_reg\[23\] GCDdpath0.B_reg\[22\] GCDdpath0.B_reg\[21\] _0536_ VGND
+ VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or4_1
X_4225_ net277 _2135_ _2129_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4156_ _2084_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3107_ _1156_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__or2_1
X_4087_ _0627_ _2018_ _0626_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__o21a_1
X_3038_ GCDdpath0.B_reg\[109\] net270 VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__or2b_1
XFILLER_0_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4989_ clknet_leaf_24_clk _0321_ _0065_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 operands_bits_A[112] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 operands_bits_A[122] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput37 operands_bits_A[17] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
Xinput48 operands_bits_A[27] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_107_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput59 operands_bits_A[37] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4010_ net45 _1957_ _1898_ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4912_ _2460_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4843_ _2449_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4774_ _2438_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3725_ net90 _1414_ _1508_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3656_ GCDdpath0.B_reg\[75\] _1654_ _1442_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ _0656_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or2b_1
XFILLER_0_141_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3587_ _0900_ _0906_ _1574_ _1576_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_73_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2538_ net365 GCDdpath0.B_reg\[7\] VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2469_ GCDdpath0.B_reg\[63\] GCDdpath0.B_reg\[62\] GCDdpath0.B_reg\[61\] GCDdpath0.B_reg\[60\]
+ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or4_1
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4208_ net283 _2123_ _2115_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__mux2_1
X_4139_ _2064_ _2069_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3510_ _1014_ _1528_ _0858_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4490_ net318 _2322_ _2316_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3441_ net6 _1467_ _1468_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3372_ _1407_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__clkbuf_4
X_5111_ clknet_leaf_38_clk _0443_ _0187_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ clknet_leaf_5_clk _0374_ _0118_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4826_ _2446_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4757_ _2435_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3708_ _0947_ _0946_ _1675_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4688_ _2424_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3639_ net104 _1640_ _1565_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput205 operands_bits_B[53] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
Xinput216 operands_bits_B[63] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
Xinput227 operands_bits_B[73] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_1
Xinput238 operands_bits_B[83] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_145_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 operands_bits_B[93] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_162_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 net325 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3990_ _0639_ _0640_ _0703_ _1940_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__nor4_1
XFILLER_0_174_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2941_ _0931_ _0938_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__or3_1
XFILLER_0_174_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2872_ _0919_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4611_ net396 _2406_ _2044_ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4542_ _2359_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4473_ _2310_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3424_ _1021_ _1453_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3355_ _1292_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__buf_2
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3286_ net27 _1305_ _1306_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__o21a_1
X_5025_ clknet_leaf_9_clk _0357_ _0101_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4809_ _2444_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_168_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ _1187_ _1190_ _0727_ _0725_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3071_ _1093_ _1121_ _1094_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_173_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3973_ net52 _1804_ _0516_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2924_ _0946_ _0950_ _0957_ _0974_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__nor4_1
XFILLER_0_85_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2855_ _0905_ GCDdpath0.B_reg\[82\] VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__nor2_2
XFILLER_0_171_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2786_ _0823_ _0826_ _0832_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__and4_2
XFILLER_0_115_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4525_ _2347_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4456_ _2298_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3407_ net11 _1341_ _1342_ _1439_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__o31a_1
X_4387_ _0564_ net220 _2242_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3338_ _1103_ _1373_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_142_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _1148_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5008_ clknet_leaf_24_clk _0340_ _0084_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_163_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2640_ GCDdpath0.B_reg\[22\] VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2571_ _0620_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput306 net306 VGND VGND VPWR VPWR result_bits_data[26] sky130_fd_sc_hd__clkbuf_4
Xoutput317 net317 VGND VGND VPWR VPWR result_bits_data[36] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput328 net328 VGND VGND VPWR VPWR result_bits_data[46] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4310_ net377 _2195_ _2187_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput339 net339 VGND VGND VPWR VPWR result_bits_data[56] sky130_fd_sc_hd__buf_2
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4241_ _2147_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4172_ net51 _1496_ _1508_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__a21o_1
X_3123_ _0624_ _0638_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3054_ net281 GCDdpath0.B_reg\[119\] VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3956_ net313 _1910_ _1911_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2907_ net355 GCDdpath0.B_reg\[70\] VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3887_ _0786_ _1848_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2838_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2769_ GCDdpath0.B_reg\[34\] net315 VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4508_ _2335_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4439_ _2272_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3810_ net336 _1539_ _1786_ _1306_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4790_ _2441_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_18 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _0722_ _1727_ _0720_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3672_ _0941_ _0986_ _1627_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_97_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2623_ net298 GCDdpath0.B_reg\[19\] VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_11_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2554_ net293 GCDdpath0.B_reg\[14\] VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_58_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2485_ GCDdpath0.B_reg\[20\] VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4224_ GCDdpath0.B_reg\[115\] net146 _2127_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4155_ _2079_ _2083_ _1288_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__mux2_1
X_3106_ net290 _1155_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4086_ _2024_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3037_ _1082_ _1040_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4988_ clknet_leaf_23_clk _0320_ _0064_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3939_ GCDdpath0.B_reg\[34\] _1896_ _1892_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput16 operands_bits_A[113] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 operands_bits_A[123] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput38 operands_bits_A[18] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_1
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput49 operands_bits_A[28] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
XFILLER_0_123_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4911_ _2460_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4842_ _2449_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4773_ _2438_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3724_ GCDdpath0.B_reg\[65\] _1409_ _1712_ _1412_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3655_ _0915_ _1653_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2606_ net308 GCDdpath0.B_reg\[28\] VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3586_ net112 _1341_ _1342_ _1594_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__o31a_1
XFILLER_0_141_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2537_ GCDdpath0.B_reg\[7\] net365 VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2468_ GCDdpath0.B_reg\[59\] GCDdpath0.B_reg\[58\] GCDdpath0.B_reg\[57\] GCDdpath0.B_reg\[56\]
+ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or4_1
X_4207_ GCDdpath0.B_reg\[120\] net152 _2113_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__mux2_1
X_4138_ _0602_ GCDdpath0.B_reg\[6\] _2068_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4069_ _1764_ _1962_ _2007_ _2008_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_137_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ _1336_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__buf_2
XFILLER_0_123_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3371_ _1302_ _1406_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5110_ clknet_leaf_25_clk _0442_ _0186_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_155_Left_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5041_ clknet_leaf_5_clk _0373_ _0117_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4825_ _2446_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4756_ _2435_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_3707_ _1698_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4687_ _2424_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3638_ GCDdpath0.B_reg\[78\] _1639_ _1598_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3569_ _0886_ _1579_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput206 operands_bits_B[54] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
Xinput217 operands_bits_B[64] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
Xinput228 operands_bits_B[74] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__buf_1
Xinput239 operands_bits_B[84] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_145_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 GCDdpath0.B_reg\[9\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2940_ _0914_ _0917_ _0989_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__o211a_1
XFILLER_0_168_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2871_ _0920_ _0921_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4610_ GCDdpath0.B_reg\[0\] net129 _1495_ VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4541_ net302 _2357_ _2358_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4472_ net324 _2309_ _2301_ VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3423_ _1084_ _1447_ _1250_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3354_ net17 _1391_ _1337_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3285_ GCDdpath0.B_reg\[123\] _1325_ _1327_ _1331_ _1303_ VGND VGND VPWR VPWR _1332_
+ sky130_fd_sc_hd__o221a_1
X_5024_ clknet_leaf_10_clk _0356_ _0100_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_135_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4808_ _2440_ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4739_ _2432_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3070_ GCDdpath0.B_reg\[114\] net276 VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__and2b_1
XFILLER_0_173_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3972_ GCDdpath0.B_reg\[30\] _1925_ _1797_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2923_ _0965_ _0969_ _0973_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2854_ net368 VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2785_ _0834_ _0835_ _0779_ _0792_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4524_ net307 _2346_ _2344_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4455_ net329 _2297_ _2287_ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3406_ net270 _1293_ _1438_ _1308_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4386_ _2249_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3337_ net279 _1324_ _1376_ _1377_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_142_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _1141_ _1144_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ clknet_leaf_15_clk _0339_ _0083_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_3199_ net266 GCDdpath0.B_reg\[105\] VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_83_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_101_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_110_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2570_ net271 GCDdpath0.B_reg\[10\] VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput307 net307 VGND VGND VPWR VPWR result_bits_data[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput318 net318 VGND VGND VPWR VPWR result_bits_data[37] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput329 net329 VGND VGND VPWR VPWR result_bits_data[47] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4240_ net273 _2146_ _2144_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4171_ GCDdpath0.B_reg\[2\] _1327_ _2096_ _1412_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__a211o_1
X_3122_ _0697_ _0649_ _1172_ _0647_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3053_ _1099_ _1100_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3955_ _1601_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__buf_2
XFILLER_0_86_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2906_ _0953_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3886_ net325 _1793_ _1851_ _0573_ _1852_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2837_ _0886_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2768_ GCDdpath0.B_reg\[35\] net316 VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4507_ net313 _2334_ _2330_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__mux2_1
X_2699_ _0748_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_76_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4438_ GCDdpath0.B_reg\[52\] net204 _2285_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4369_ _2237_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3740_ _0838_ _1726_ _0728_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3671_ _1667_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2622_ net297 GCDdpath0.B_reg\[18\] VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2553_ _0588_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_58_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2484_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or3_1
X_4223_ _2134_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4154_ GCDdpath0.B_reg\[5\] _2081_ _2082_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3105_ net290 _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4085_ net294 _2023_ _1992_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3036_ _1017_ _1083_ _1085_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4987_ clknet_leaf_23_clk _0319_ _0063_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3938_ _0761_ _1889_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3869_ _0778_ _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_115_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 operands_bits_A[114] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 operands_bits_A[124] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_0_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput39 operands_bits_A[19] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_109_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4910_ _2460_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4841_ _2449_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4772_ _2433_ VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3723_ _1549_ _1711_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3654_ _0916_ _1222_ _1652_ _1223_ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2605_ GCDdpath0.B_reg\[28\] net308 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3585_ net371 _1539_ _1593_ _1308_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2536_ net321 GCDdpath0.B_reg\[3\] VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2467_ GCDctrl0.state\[1\] VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__inv_2
X_4206_ _2122_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4137_ _0590_ _2067_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4068_ GCDdpath0.B_reg\[16\] _1520_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3019_ _1043_ _1069_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3370_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_90_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5040_ clknet_leaf_6_clk _0372_ _0116_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4824_ _2446_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4755_ _2435_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3706_ net352 _1697_ _1687_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4686_ _2419_ VGND VGND VPWR VPWR _2424_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3637_ _0937_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3568_ _0885_ _1577_ _0889_ _1578_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_149_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2519_ _0518_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__or2_1
X_3499_ _1053_ _1421_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__or2_1
Xinput207 operands_bits_B[55] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_2
XFILLER_0_110_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput218 operands_bits_B[65] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
Xinput229 operands_bits_B[75] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_1
X_5169_ clknet_leaf_6_clk _0501_ _0245_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_162_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_162_Right_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 net278 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_162_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2870_ GCDdpath0.B_reg\[73\] net358 VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__and2b_1
XFILLER_0_127_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4540_ _1295_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4471_ GCDdpath0.B_reg\[42\] net193 _2299_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3422_ net268 _1445_ _1451_ _1452_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3353_ GCDdpath0.B_reg\[114\] _1390_ _1319_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3284_ _1130_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__xnor2_1
X_5023_ clknet_leaf_9_clk _0355_ _0099_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ _2443_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2999_ GCDdpath0.B_reg\[97\] net384 VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4738_ _2432_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4669_ _2421_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_174_Left_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_168_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3971_ _0651_ _1924_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2922_ _0970_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2853_ _0902_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2784_ _0794_ _0797_ _0793_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_171_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4523_ GCDdpath0.B_reg\[27\] net176 _2342_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4454_ GCDdpath0.B_reg\[47\] net198 _2285_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3405_ _1435_ _1436_ _1437_ GCDdpath0.B_reg\[109\] VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_141_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4385_ net352 _2248_ _2244_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3336_ net20 _1305_ _1369_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_142_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _1309_ _1315_ _1294_ net288 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_1_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ clknet_leaf_15_clk _0338_ _0082_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_3198_ _1043_ _1056_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput308 net308 VGND VGND VPWR VPWR result_bits_data[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput319 net319 VGND VGND VPWR VPWR result_bits_data[38] sky130_fd_sc_hd__buf_2
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4170_ _0585_ _1620_ _2095_ VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__and3_1
X_3121_ _0657_ _0660_ _1171_ _0659_ _0698_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__a311o_1
XFILLER_0_172_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3052_ _1101_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3954_ net54 _1909_ _1898_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2905_ _0954_ _0955_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3885_ net66 _1804_ _1734_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__or3_1
XFILLER_0_156_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2836_ net372 GCDdpath0.B_reg\[86\] VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2767_ _0762_ _0767_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_152_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4506_ GCDdpath0.B_reg\[32\] net182 _2328_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2698_ net337 GCDdpath0.B_reg\[54\] VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4437_ _2227_ VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4368_ net358 _2236_ _2230_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3319_ _1105_ _1106_ _1108_ _1361_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__or4_1
X_4299_ _2188_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3670_ net358 _1666_ _1602_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2621_ _0664_ _0667_ _0668_ _0671_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_97_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2552_ _0602_ GCDdpath0.B_reg\[6\] _0589_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2483_ GCDdpath0.B_reg\[3\] GCDdpath0.B_reg\[2\] GCDdpath0.B_reg\[1\] GCDdpath0.B_reg\[0\]
+ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4222_ net400 _2133_ _2129_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__mux2_1
X_4153_ _1319_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_71_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3104_ GCDdpath0.B_reg\[127\] VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__inv_2
X_4084_ net35 _2022_ _1984_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3035_ GCDdpath0.B_reg\[107\] net268 VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__or2b_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4986_ clknet_leaf_25_clk _0318_ _0062_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3937_ _1895_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3868_ _0773_ _1825_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2819_ _0865_ _0869_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3799_ GCDdpath0.B_reg\[55\] _1285_ _1549_ _1777_ _1340_ VGND VGND VPWR VPWR _1778_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 operands_bits_A[115] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xinput29 operands_bits_A[125] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4840_ _2449_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4771_ _2437_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3722_ _0953_ _1710_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3653_ _0988_ _1628_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2604_ _0653_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3584_ GCDdpath0.B_reg\[85\] _1437_ _1343_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__o22a_1
XFILLER_0_141_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2535_ GCDdpath0.B_reg\[3\] net321 VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_110_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2466_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4205_ net284 _2121_ _2115_ VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4136_ _0600_ _2066_ _0593_ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4067_ _1961_ _1174_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3018_ _1054_ _1061_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__or3_1
XFILLER_0_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4969_ clknet_leaf_28_clk _0301_ _0045_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4823_ _2446_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4754_ _2435_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_172_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_173_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3705_ net93 _1696_ _1665_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4685_ _2423_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3636_ _0924_ _1636_ _1630_ _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3567_ _0880_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2518_ _0543_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3498_ _1509_ _1510_ _1515_ _1518_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__o22a_1
Xinput208 operands_bits_B[56] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
Xinput219 operands_bits_B[66] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_87_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5168_ clknet_leaf_6_clk _0500_ _0244_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_166_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4119_ net271 _2052_ _2041_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__mux2_1
X_5099_ clknet_leaf_38_clk _0431_ _0175_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_123_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_764 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4470_ _2308_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3421_ net9 _1432_ _1369_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3352_ _1097_ _1383_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3283_ _1131_ _1329_ _1132_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__a21bo_1
X_5022_ clknet_leaf_10_clk _0354_ _0098_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_144_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4806_ _2443_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2998_ net384 GCDdpath0.B_reg\[97\] VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4737_ _2432_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4668_ _2421_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3619_ _0898_ _0998_ _1526_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__and3_1
X_4599_ net332 _2398_ _2044_ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_165_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3970_ _0660_ _1918_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2921_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_100_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2852_ GCDdpath0.B_reg\[81\] net367 VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ _0795_ _0798_ _0800_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__or4b_1
XFILLER_0_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4522_ _2345_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4453_ _2296_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3404_ _1284_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__buf_2
X_4384_ GCDdpath0.B_reg\[68\] net221 _2242_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3335_ GCDdpath0.B_reg\[117\] _1325_ _1327_ _1375_ _1303_ VGND VGND VPWR VPWR _1376_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_142_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3266_ _1282_ _1311_ _1312_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a31o_1
X_5005_ clknet_leaf_15_clk _0337_ _0081_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _1058_ _1065_ _1246_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_523 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput309 net309 VGND VGND VPWR VPWR result_bits_data[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_168_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3120_ _1168_ _1170_ _0640_ _0656_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3051_ GCDdpath0.B_reg\[116\] net278 VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3953_ _1464_ _1888_ _1907_ _1908_ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2904_ net348 GCDdpath0.B_reg\[64\] VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3884_ GCDdpath0.B_reg\[43\] _1850_ _1797_ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2835_ GCDdpath0.B_reg\[86\] net372 VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2766_ _0763_ _0766_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4505_ _2333_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
X_2697_ GCDdpath0.B_reg\[54\] net337 VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__and2b_1
X_4436_ _2284_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4367_ GCDdpath0.B_reg\[73\] net227 _2228_ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3318_ _1125_ _1360_ _1109_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__a21oi_1
X_4298_ net381 _2185_ _2187_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__mux2_1
X_3249_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2620_ _0669_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_97_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2551_ net354 VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2482_ GCDdpath0.B_reg\[15\] GCDdpath0.B_reg\[14\] GCDdpath0.B_reg\[13\] GCDdpath0.B_reg\[12\]
+ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_75_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4221_ GCDdpath0.B_reg\[116\] net147 _2127_ VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4152_ _0594_ _2080_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_50_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3103_ _0577_ _1150_ _1151_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4083_ GCDdpath0.B_reg\[15\] _2021_ _1989_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__mux2_1
X_3034_ _1024_ _1022_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4985_ clknet_leaf_26_clk _0317_ _0061_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3936_ net316 _1894_ _1841_ VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3867_ _1836_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2818_ _0867_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3798_ _0747_ _1776_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2749_ net318 GCDdpath0.B_reg\[37\] VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4419_ _2272_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 operands_bits_A[116] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XFILLER_0_150_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_116_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4770_ _2437_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3721_ _0954_ _1674_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3652_ _1651_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2603_ GCDdpath0.B_reg\[24\] net304 VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3583_ _1590_ _1591_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2534_ _0579_ _0582_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2465_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__clkbuf_2
X_4204_ GCDdpath0.B_reg\[121\] net153 _2113_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__mux2_1
X_4135_ _0597_ _2065_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4066_ _2006_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3017_ _1064_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4968_ clknet_leaf_36_clk _0300_ _0044_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3919_ _0801_ _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4899_ _2458_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4822_ _2440_ VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_66_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_172_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4753_ _2435_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3704_ _1280_ _1676_ _1694_ _1695_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4684_ _2423_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3635_ _0925_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3566_ _0900_ _0906_ _1574_ _1575_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__o311a_1
XFILLER_0_141_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2517_ _0556_ _0557_ _0561_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__or4_2
X_3497_ GCDdpath0.B_reg\[97\] _1516_ _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput209 operands_bits_B[57] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
X_5167_ clknet_leaf_3_clk _0499_ _0243_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_162_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4118_ net12 _2051_ _2029_ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__mux2_1
X_5098_ clknet_2_1__leaf_clk _0430_ _0174_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4049_ _1601_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_123_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3420_ GCDdpath0.B_reg\[107\] _1417_ _1418_ _1450_ _1387_ VGND VGND VPWR VPWR _1451_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3351_ net277 _1324_ _1388_ _1389_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3282_ _1142_ _1328_ _1135_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a21oi_1
X_5021_ clknet_leaf_10_clk _0353_ _0097_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_144_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4805_ _2443_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2997_ _1046_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4736_ _2426_ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4667_ _2421_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3618_ _1622_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_1
X_4598_ GCDdpath0.B_reg\[4\] net201 _1495_ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3549_ _0875_ _0871_ _0873_ _1551_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_164_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2920_ GCDdpath0.B_reg\[68\] net352 VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__or2b_1
XFILLER_0_168_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2851_ net367 GCDdpath0.B_reg\[81\] VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2782_ _0799_ _0802_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ net308 _2343_ _2344_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4452_ net330 _2295_ _2287_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3403_ _1036_ _1082_ _1434_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4383_ _2247_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3334_ _1371_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__xnor2_1
X_3265_ GCDdpath0.B_reg\[125\] _1313_ _1288_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5004_ clknet_leaf_18_clk _0336_ _0080_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_3196_ _1057_ _1059_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4719_ _2429_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3050_ net278 GCDdpath0.B_reg\[116\] VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__and2b_1
XFILLER_0_171_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3952_ GCDdpath0.B_reg\[32\] _1464_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2903_ GCDdpath0.B_reg\[64\] net348 VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3883_ _0782_ _1849_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2834_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2765_ _0746_ _0809_ _0751_ _0814_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4504_ net314 _2332_ _2330_ VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2696_ _0745_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4435_ net336 _2283_ _2273_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4366_ _2235_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3317_ _1122_ _1359_ _1104_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__a21o_1
X_4297_ _2186_ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__buf_2
X_3248_ _0518_ _1284_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__nor2_1
X_3179_ _0896_ _1004_ _0903_ _0906_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2550_ _0591_ _0593_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2481_ GCDdpath0.B_reg\[11\] GCDdpath0.B_reg\[10\] GCDdpath0.B_reg\[9\] GCDdpath0.B_reg\[8\]
+ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4220_ _2132_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_1
X_4151_ _0595_ _2066_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3102_ _0575_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4082_ _0606_ _2020_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__xor2_1
X_3033_ _1023_ _1025_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4984_ clknet_leaf_38_clk _0316_ _0060_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3935_ net57 _1893_ _1817_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3866_ _1831_ _1835_ _1340_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2817_ _0866_ GCDdpath0.B_reg\[90\] VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3797_ _0749_ _1775_ _0809_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2748_ GCDdpath0.B_reg\[37\] net318 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2679_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4418_ _1395_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4349_ GCDdpath0.B_reg\[78\] net232 _2213_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3720_ _1709_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3651_ net361 _1650_ _1602_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2602_ net304 GCDdpath0.B_reg\[24\] VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3582_ _0883_ _1577_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2533_ _0578_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ net257 net259 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nand2_2
XFILLER_0_139_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4203_ _2120_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4134_ _0578_ _0585_ _0586_ _0587_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4065_ net296 _2005_ _1992_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3016_ _1065_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_125_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4967_ clknet_leaf_31_clk _0299_ _0043_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3918_ _0802_ _1869_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_163_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4898_ _2458_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3849_ net329 net70 _1496_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_172_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_167_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4821_ _2445_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4752_ _2435_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3703_ GCDdpath0.B_reg\[68\] _1520_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__and2_1
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4683_ _2423_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3634_ GCDdpath0.B_reg\[76\] net361 VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3565_ net369 GCDdpath0.B_reg\[83\] VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2516_ _0562_ _0563_ _0565_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_149_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3496_ _0572_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__buf_2
XFILLER_0_166_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5166_ clknet_leaf_7_clk _0498_ _0242_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_127_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4117_ _1764_ _2016_ _2049_ _2050_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_162_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5097_ clknet_leaf_30_clk _0429_ _0173_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dfrtp_4
X_4048_ net39 _1990_ _1984_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_169_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput290 net290 VGND VGND VPWR VPWR result_bits_data[127] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_167_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3350_ net18 _1305_ _1369_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3281_ _1118_ _1127_ _1139_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a21o_1
X_5020_ clknet_leaf_10_clk _0352_ _0096_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4804_ _2443_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2996_ net385 GCDdpath0.B_reg\[98\] VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__xor2_2
XFILLER_0_174_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4735_ _2431_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4666_ _2421_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
X_3617_ _1616_ _1621_ _1340_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4597_ _2397_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3548_ _0875_ _0871_ _0873_ _1551_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_164_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3479_ _1046_ _1501_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_134_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5149_ clknet_leaf_12_clk _0481_ _0225_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_143_Left_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Left_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_161_Left_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2850_ _0899_ _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2781_ _0827_ _0526_ _0828_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__o31a_1
X_4520_ _2272_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__buf_2
XFILLER_0_170_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4451_ GCDdpath0.B_reg\[48\] net199 _2285_ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_170_Left_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3402_ _1036_ _1082_ _1434_ _1280_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__o31a_1
X_4382_ net353 _2246_ _2244_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3333_ _1372_ _1373_ _1102_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3264_ _1284_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5003_ clknet_leaf_18_clk _0335_ _0079_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3195_ _1062_ _1245_ _1066_ _1063_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2979_ net273 GCDdpath0.B_reg\[111\] VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4718_ _2429_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4649_ _2417_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3951_ _0765_ _0684_ _0708_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2902_ _0951_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3882_ _0785_ _0786_ _1848_ _0784_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__o31a_1
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2833_ _0882_ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_170_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2764_ _0745_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4503_ GCDdpath0.B_reg\[33\] net183 _2328_ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2695_ net338 GCDdpath0.B_reg\[55\] VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__and2b_1
X_4434_ GCDdpath0.B_reg\[53\] net205 _2270_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4365_ net359 _2234_ _2230_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_171_Right_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3316_ _1120_ _1358_ _1098_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4296_ _1395_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__buf_2
X_3247_ _1153_ _0577_ _1150_ _1151_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__or4_1
XFILLER_0_174_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3178_ _0880_ _0881_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2480_ GCDdpath0.B_reg\[7\] GCDdpath0.B_reg\[6\] GCDdpath0.B_reg\[5\] GCDdpath0.B_reg\[4\]
+ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_75_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4150_ net343 net84 _1615_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3101_ net289 GCDdpath0.B_reg\[126\] VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__and2b_1
X_4081_ net293 _2012_ _2019_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3032_ GCDdpath0.B_reg\[106\] net267 VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__or2b_1
Xinput190 operands_bits_B[3] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4983_ clknet_leaf_38_clk _0315_ _0059_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3934_ GCDdpath0.B_reg\[35\] _1891_ _1892_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3865_ _0526_ _1833_ _1834_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_171_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2816_ _0866_ GCDdpath0.B_reg\[90\] VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3796_ _0813_ _1774_ _0752_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_115_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2747_ _0796_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_132_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2678_ _0725_ _0726_ _0727_ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__and4_1
XFILLER_0_140_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4417_ GCDdpath0.B_reg\[58\] net210 _2270_ VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4348_ _2222_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_1
X_4279_ GCDdpath0.B_reg\[99\] net255 _2170_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3650_ net102 _1649_ _1565_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2601_ _0647_ _0648_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_77_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3581_ _0880_ _0882_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2532_ net310 GCDdpath0.B_reg\[2\] VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2463_ _2409_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__inv_2
X_4202_ net285 _2119_ _2115_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5182_ clknet_leaf_26_clk _0514_ _0258_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4133_ _0588_ _0589_ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_147_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4064_ net37 _2004_ _1984_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3015_ net262 GCDdpath0.B_reg\[101\] VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__or2b_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4966_ clknet_leaf_31_clk _0298_ _0042_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3917_ net318 net59 _1615_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4897_ _2458_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3848_ _1819_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3779_ _0713_ _1747_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__and2b_1
XFILLER_0_171_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4820_ _2445_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4751_ _2433_ VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3702_ _0973_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4682_ _2423_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3633_ net364 _1349_ _1634_ _1635_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3564_ _0881_ _0883_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2515_ GCDdpath0.B_reg\[71\] GCDdpath0.B_reg\[70\] GCDdpath0.B_reg\[69\] GCDdpath0.B_reg\[68\]
+ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_149_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3495_ _1300_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__clkbuf_4
X_5165_ clknet_leaf_3_clk _0497_ _0241_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_166_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4116_ GCDdpath0.B_reg\[10\] _1398_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_162_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5096_ clknet_leaf_36_clk _0428_ _0172_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_162_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4047_ GCDdpath0.B_reg\[19\] _1988_ _1989_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4949_ clknet_leaf_43_clk _0281_ _0025_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_164_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_65_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput280 net280 VGND VGND VPWR VPWR result_bits_data[118] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput291 net291 VGND VGND VPWR VPWR result_bits_data[12] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_167_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3280_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_144_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4803_ _2443_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2995_ _1044_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4734_ _2431_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4665_ _2419_ VGND VGND VPWR VPWR _2421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3616_ _1618_ _1619_ _1620_ GCDdpath0.B_reg\[81\] VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_102_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4596_ net343 _2396_ _2386_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3547_ net377 _1440_ _1558_ _1559_ _1560_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__o221a_1
XFILLER_0_101_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3478_ _1072_ _0553_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5148_ clknet_leaf_12_clk _0480_ _0224_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_4_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5079_ clknet_leaf_41_clk _0411_ _0155_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_167_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2780_ _0772_ _0829_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_143_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4450_ _2294_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__clkbuf_1
X_3401_ _1041_ _1423_ _1040_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__o21ai_1
X_4381_ GCDdpath0.B_reg\[69\] net222 _2242_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3332_ _1122_ _1359_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3263_ _0577_ _1145_ _1147_ _1310_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_147_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5002_ clknet_leaf_20_clk _0334_ _0078_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
X_3194_ net385 _1242_ _1244_ _1044_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2978_ GCDdpath0.B_reg\[111\] net273 VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4717_ _2429_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4648_ _2417_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4579_ GCDdpath0.B_reg\[10\] net140 _2384_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_165_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3950_ _1906_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2901_ GCDdpath0.B_reg\[65\] net349 VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__and2b_1
XFILLER_0_129_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3881_ _0791_ _1823_ _0787_ _0790_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2832_ GCDdpath0.B_reg\[84\] net370 VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2763_ _0757_ _0811_ _0812_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4502_ _2331_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2694_ GCDdpath0.B_reg\[55\] net338 VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_152_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4433_ _2282_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4364_ GCDdpath0.B_reg\[74\] net228 _2228_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3315_ _1071_ _1092_ _1112_ _1115_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__a211o_1
X_4295_ GCDdpath0.B_reg\[94\] net250 _2184_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__mux2_1
X_3246_ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3177_ _0942_ _0963_ _1219_ _1227_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_174_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3100_ _1145_ _1147_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4080_ _0627_ _2018_ _0605_ _0626_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__o211a_1
X_3031_ _1037_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__clkbuf_2
Xinput180 operands_bits_B[30] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_1
XFILLER_0_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput191 operands_bits_B[40] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_1
XFILLER_0_163_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4982_ clknet_leaf_25_clk _0314_ _0058_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3933_ _1318_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3864_ _1279_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2815_ net377 VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3795_ _0755_ _1773_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_115_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2746_ GCDdpath0.B_reg\[38\] net319 VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2677_ GCDdpath0.B_reg\[61\] net345 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4416_ _2227_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4347_ net364 _2221_ _2215_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__mux2_1
X_4278_ _2173_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3229_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2600_ _0649_ _0650_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3580_ net372 _1349_ _1588_ _1589_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2531_ net394 _0580_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2462_ _2409_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4201_ GCDdpath0.B_reg\[122\] net154 _2113_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5181_ clknet_leaf_13_clk _0513_ _0257_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4132_ _2063_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4063_ GCDdpath0.B_reg\[17\] _2003_ _1989_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3014_ GCDdpath0.B_reg\[101\] net262 VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_108_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4965_ clknet_leaf_31_clk _0297_ _0041_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3916_ net319 _1793_ _1876_ _0573_ _1877_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4896_ _2458_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3847_ net330 _1818_ _1745_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_171_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3778_ net340 net81 _1496_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2729_ net325 GCDdpath0.B_reg\[43\] VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4750_ _2434_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3701_ _0978_ _1675_ _0944_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4681_ _2423_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3632_ net105 _1583_ _1517_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_153_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3563_ _1006_ _1573_ _1004_ _0909_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2514_ _0564_ GCDdpath0.B_reg\[66\] GCDdpath0.B_reg\[65\] GCDdpath0.B_reg\[64\] VGND
+ VGND VPWR VPWR _0565_ sky130_fd_sc_hd__or4_1
X_3494_ _1511_ _1514_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_149_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5164_ clknet_leaf_3_clk _0496_ _0240_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_166_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4115_ _0621_ _2015_ VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5095_ clknet_leaf_30_clk _0427_ _0171_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_162_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4046_ _1278_ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_166_Right_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4948_ clknet_leaf_40_clk _0280_ _0024_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4879_ _2455_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput270 net270 VGND VGND VPWR VPWR result_bits_data[109] sky130_fd_sc_hd__clkbuf_4
Xoutput281 net281 VGND VGND VPWR VPWR result_bits_data[119] sky130_fd_sc_hd__clkbuf_4
Xoutput292 net292 VGND VGND VPWR VPWR result_bits_data[13] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4802_ _2443_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2994_ GCDdpath0.B_reg\[99\] net386 VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__or2b_1
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4733_ _2431_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4664_ _2420_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3615_ _1395_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4595_ GCDdpath0.B_reg\[5\] net212 _2384_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3546_ net118 _1506_ _1355_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3477_ _1047_ _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_164_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5147_ clknet_leaf_10_clk _0479_ _0223_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_4_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5078_ clknet_leaf_41_clk _0410_ _0154_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4029_ GCDdpath0.B_reg\[22\] _1409_ _1974_ _1412_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3400_ net272 _1324_ _1431_ _1433_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4380_ _2245_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3331_ _1101_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_84_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3262_ _0577_ _1145_ _1147_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5001_ clknet_leaf_20_clk _0333_ _0077_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3193_ _1048_ _1050_ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_93_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2977_ _1022_ _1023_ _1024_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_174_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4716_ _2429_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4647_ _2417_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4578_ _2313_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3529_ _1529_ _1544_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_164_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2900_ net349 GCDdpath0.B_reg\[65\] VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__and2b_2
XFILLER_0_168_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3880_ net67 _1354_ _1414_ _1847_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2831_ GCDdpath0.B_reg\[85\] net371 VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__and2b_1
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2762_ GCDdpath0.B_reg\[53\] net336 VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4501_ net315 _2329_ _2330_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2693_ _0741_ _0742_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4432_ net337 _2281_ _2273_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4363_ _2233_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3314_ net22 _0517_ _1308_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4294_ _2141_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3245_ _1279_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__buf_2
X_3176_ _0993_ _0936_ _1226_ _0932_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__a31o_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_802 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Left_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_158_Left_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3030_ _1029_ _1031_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__and2b_1
Xinput170 operands_bits_B[21] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xinput181 operands_bits_B[31] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
Xinput192 operands_bits_B[41] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4981_ clknet_leaf_27_clk _0313_ _0057_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_3932_ _0760_ _1890_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3863_ _0771_ _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Left_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2814_ _0863_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3794_ _0810_ _1772_ _0742_ _0756_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2745_ net319 GCDdpath0.B_reg\[38\] VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__and2b_1
XFILLER_0_147_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2676_ net345 GCDdpath0.B_reg\[61\] VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4415_ _2269_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4346_ GCDdpath0.B_reg\[79\] net233 _2213_ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__mux2_1
X_4277_ net261 _2171_ _2172_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__mux2_1
X_3228_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_154_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3159_ _1206_ _1207_ _1209_ _0759_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2530_ net299 GCDdpath0.B_reg\[1\] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4200_ _2118_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__clkbuf_1
X_5180_ clknet_leaf_13_clk _0512_ _0256_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4131_ net376 _2062_ _2041_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4062_ _2001_ _2002_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3013_ _1062_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_108_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4964_ clknet_leaf_32_clk _0296_ _0040_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3915_ net60 _1804_ _1734_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4895_ _2458_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3846_ net71 _1816_ _1817_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3777_ _1758_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_171_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2728_ _0772_ _0775_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__or3_2
XFILLER_0_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2659_ net392 GCDdpath0.B_reg\[58\] VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4329_ GCDdpath0.B_reg\[84\] net239 _2199_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3700_ net94 _1341_ _1342_ _1692_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4680_ _2423_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3631_ GCDdpath0.B_reg\[79\] _1285_ _1549_ _1633_ _1536_ VGND VGND VPWR VPWR _1634_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3562_ _0998_ _1526_ _0898_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2513_ GCDdpath0.B_reg\[67\] VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3493_ _1512_ _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_149_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_166_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5163_ clknet_leaf_12_clk _0495_ _0239_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dfrtp_4
X_4114_ _1509_ _2043_ _2047_ _2048_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5094_ clknet_leaf_30_clk _0426_ _0170_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_127_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4045_ _0674_ _1987_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ clknet_leaf_42_clk _0279_ _0023_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4878_ _2455_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3829_ GCDdpath0.B_reg\[50\] _1802_ _1797_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_171_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_719 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput260 net394 VGND VGND VPWR VPWR result_bits_data[0] sky130_fd_sc_hd__clkbuf_4
Xoutput271 net271 VGND VGND VPWR VPWR result_bits_data[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput282 net282 VGND VGND VPWR VPWR result_bits_data[11] sky130_fd_sc_hd__clkbuf_4
Xoutput293 net293 VGND VGND VPWR VPWR result_bits_data[14] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4801_ _2440_ VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2993_ net386 GCDdpath0.B_reg\[99\] VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4732_ _2431_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4663_ _2420_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3614_ _0904_ _1617_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4594_ _2395_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3545_ _1353_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__clkbuf_4
X_3476_ _1074_ _1498_ _1049_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_164_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5146_ clknet_leaf_12_clk _0478_ _0222_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5077_ clknet_leaf_40_clk _0409_ _0153_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dfrtp_1
X_4028_ _1620_ _1966_ _1973_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__and3_1
XFILLER_0_67_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3330_ _1099_ _1100_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3261_ _1141_ _1144_ _1148_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__a21oi_1
X_5000_ clknet_leaf_20_clk _0332_ _0076_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3192_ _1051_ _1049_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2976_ _1025_ _1026_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4715_ _2426_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4646_ _2417_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4577_ _2383_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3528_ _0858_ _1014_ _1528_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__and3_1
X_3459_ net263 _1484_ _1393_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__mux2_1
X_5129_ clknet_leaf_20_clk _0461_ _0205_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_164_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2830_ net370 GCDdpath0.B_reg\[84\] VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__and2b_1
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2761_ _0752_ _0755_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__or2b_1
XFILLER_0_27_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4500_ _2272_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2692_ GCDdpath0.B_reg\[51\] net334 VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_1 operands_bits_B[50] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4431_ GCDdpath0.B_reg\[54\] net206 _2270_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4362_ net360 _2232_ _2230_ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3313_ net283 _1349_ _1352_ _1354_ _1356_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _2183_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__clkbuf_1
X_3244_ _0574_ _1290_ _1294_ net290 VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__o2bb2a_1
X_3175_ _0925_ _1220_ _1225_ _0935_ _0994_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_159_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2959_ GCDdpath0.B_reg\[86\] _0890_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4629_ _2413_ VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput160 operands_bits_B[12] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput171 operands_bits_B[22] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
Xinput182 operands_bits_B[32] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_1
Xinput193 operands_bits_B[42] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
X_4980_ clknet_leaf_27_clk _0312_ _0056_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_129_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3931_ _0761_ _1889_ _0820_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3862_ _0777_ _1826_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_154_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2813_ GCDdpath0.B_reg\[91\] net378 VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_171_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3793_ _0737_ _1771_ _0741_ _0733_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2744_ _0793_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2675_ GCDdpath0.B_reg\[60\] net344 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__or2b_1
XFILLER_0_169_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4414_ net342 _2268_ _2258_ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4345_ _2220_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_1
X_4276_ _2082_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3227_ _0518_ _1277_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3158_ _0830_ _1208_ _0828_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_90_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3089_ _1134_ _1135_ _1136_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4130_ net117 _2061_ _2029_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__mux2_1
X_4061_ _0676_ _1962_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3012_ net261 GCDdpath0.B_reg\[100\] VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4963_ clknet_leaf_31_clk _0295_ _0039_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3914_ GCDdpath0.B_reg\[38\] _1875_ _1797_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4894_ _2454_ VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3845_ _1336_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3776_ net392 _1757_ _1745_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2727_ _0776_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2658_ net342 GCDdpath0.B_reg\[59\] VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2589_ GCDdpath0.B_reg\[27\] net307 VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__nor2b_2
XTAP_TAPCELL_ROW_35_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4328_ _2208_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__clkbuf_1
X_4259_ GCDdpath0.B_reg\[105\] net135 _2156_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_163_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3630_ _0934_ _1632_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3561_ _1572_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2512_ GCDdpath0.B_reg\[79\] GCDdpath0.B_reg\[78\] GCDdpath0.B_reg\[77\] GCDdpath0.B_reg\[76\]
+ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3492_ _1053_ _1421_ _1052_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5162_ clknet_leaf_7_clk _0494_ _0238_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4113_ GCDdpath0.B_reg\[11\] _1516_ _1353_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__a21o_1
X_5093_ clknet_leaf_30_clk _0425_ _0169_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_127_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4044_ _0686_ _1963_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4946_ clknet_leaf_42_clk _0278_ _0022_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_163_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4877_ _2455_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3828_ _1772_ _1801_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3759_ GCDdpath0.B_reg\[60\] _1742_ _1684_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput261 net261 VGND VGND VPWR VPWR result_bits_data[100] sky130_fd_sc_hd__clkbuf_4
Xoutput272 net272 VGND VGND VPWR VPWR result_bits_data[110] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput283 net283 VGND VGND VPWR VPWR result_bits_data[120] sky130_fd_sc_hd__clkbuf_4
Xoutput294 net294 VGND VGND VPWR VPWR result_bits_data[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4800_ _2442_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2992_ _1028_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4731_ _2431_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4662_ _2420_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3613_ _0904_ _1617_ _1280_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4593_ net354 _2394_ _2386_ VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3544_ GCDdpath0.B_reg\[90\] _1557_ _1442_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3475_ _1053_ _1421_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5145_ clknet_leaf_17_clk _0477_ _0221_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_4_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5076_ clknet_leaf_40_clk _0408_ _0152_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4027_ _0664_ _1972_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4929_ clknet_leaf_40_clk _0261_ _0005_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3260_ net29 _0517_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__o21ai_1
X_3191_ _0553_ _1045_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_163_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2975_ net265 GCDdpath0.B_reg\[104\] VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__or2b_1
XFILLER_0_173_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4714_ _2428_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4645_ _2417_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4576_ net282 _2382_ _2372_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3527_ net121 _1341_ _1342_ _1543_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__o31a_1
XFILLER_0_0_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3458_ net4 _1483_ _1468_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__mux2_1
X_3389_ _1041_ _1423_ _1089_ _1040_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__o211a_1
X_5128_ clknet_leaf_21_clk _0460_ _0204_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_169_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5059_ clknet_leaf_49_clk _0391_ _0135_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2760_ _0733_ _0737_ _0744_ _0810_ _0742_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__o32a_1
XFILLER_0_143_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2691_ net334 GCDdpath0.B_reg\[51\] VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_152_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4430_ _2280_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_2 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4361_ GCDdpath0.B_reg\[75\] net229 _2228_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3312_ net24 _1288_ _1355_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_130_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4292_ net382 _2182_ _2172_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__mux2_1
X_3243_ _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3174_ _1221_ _0916_ _1224_ _0927_ _0913_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a311o_1
XFILLER_0_117_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2958_ _0880_ _0884_ _0893_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2889_ GCDdpath0.B_reg\[72\] net357 VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4628_ _2414_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4559_ GCDdpath0.B_reg\[16\] net164 _2370_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput150 operands_bits_B[119] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xinput161 operands_bits_B[13] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput172 operands_bits_B[23] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_1
Xinput183 operands_bits_B[33] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
Xinput194 operands_bits_B[43] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3930_ _0817_ _1888_ _1195_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_86_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ net328 net69 _1615_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2812_ net378 GCDdpath0.B_reg\[91\] VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3792_ _0837_ _1722_ _1770_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2743_ net320 GCDdpath0.B_reg\[39\] VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__or2b_1
XFILLER_0_125_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2674_ net344 GCDdpath0.B_reg\[60\] VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4413_ GCDdpath0.B_reg\[59\] net211 _2256_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4344_ net366 _2219_ _2215_ VGND VGND VPWR VPWR _2220_ sky130_fd_sc_hd__mux2_1
X_4275_ GCDdpath0.B_reg\[100\] net130 _2170_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3226_ _1260_ _1275_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3157_ _0827_ _0526_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3088_ _1137_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_162_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_165_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4060_ _0677_ _2000_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3011_ GCDdpath0.B_reg\[100\] net261 VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__and2b_1
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4962_ clknet_leaf_34_clk _0294_ _0038_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_114_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3913_ _0798_ _1870_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4893_ _2457_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3844_ GCDdpath0.B_reg\[48\] _1815_ _1810_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3775_ _1755_ _1756_ net82 _0571_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2726_ net327 GCDdpath0.B_reg\[45\] VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_113_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2657_ _0696_ _0699_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2588_ net307 GCDdpath0.B_reg\[27\] VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__nor2b_2
XTAP_TAPCELL_ROW_35_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4327_ net371 _2207_ _2201_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4258_ _2159_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__clkbuf_1
X_3209_ _1213_ _1256_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a21bo_1
X_4189_ _2110_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_173_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_172_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3560_ net374 _1571_ _1489_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2511_ GCDdpath0.B_reg\[75\] GCDdpath0.B_reg\[74\] GCDdpath0.B_reg\[73\] GCDdpath0.B_reg\[72\]
+ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3491_ _1049_ _1050_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5161_ clknet_leaf_6_clk _0493_ _0237_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4112_ _2044_ _2045_ _2046_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5092_ clknet_leaf_36_clk _0424_ _0168_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_127_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4043_ _1986_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4945_ clknet_leaf_44_clk _0277_ _0021_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4876_ _2455_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3827_ _0741_ _1800_ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3758_ _1741_ _1725_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2709_ net316 GCDdpath0.B_reg\[35\] VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__xor2_1
X_3689_ _0960_ _1677_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput262 net262 VGND VGND VPWR VPWR result_bits_data[101] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput273 net273 VGND VGND VPWR VPWR result_bits_data[111] sky130_fd_sc_hd__clkbuf_4
Xoutput284 net284 VGND VGND VPWR VPWR result_bits_data[121] sky130_fd_sc_hd__clkbuf_4
Xoutput295 net295 VGND VGND VPWR VPWR result_bits_data[16] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire389 _1266_ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2991_ _1035_ _1036_ _1037_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4730_ _2431_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4661_ _2420_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3612_ _1005_ _1573_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4592_ GCDdpath0.B_reg\[6\] net223 _2384_ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3543_ _0869_ _1552_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3474_ net386 net127 _1496_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5144_ clknet_leaf_17_clk _0476_ _0220_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5075_ clknet_leaf_42_clk _0407_ _0151_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dfrtp_4
X_4026_ _0694_ _1965_ _0669_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4928_ clknet_leaf_40_clk _0260_ _0004_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4859_ _2452_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _0912_ _1228_ _1237_ _0849_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_53_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_163_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2974_ GCDdpath0.B_reg\[104\] net265 VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4713_ _2428_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4644_ _2417_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4575_ GCDdpath0.B_reg\[11\] net151 _2370_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3526_ net380 _1539_ _1542_ _1308_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3457_ GCDdpath0.B_reg\[102\] _1481_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux2_1
X_3388_ _1028_ _1422_ _1087_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_71_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5127_ clknet_leaf_21_clk _0459_ _0203_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5058_ clknet_leaf_0_clk _0390_ _0134_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4009_ GCDdpath0.B_reg\[24\] _1956_ _1892_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_949 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_695 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2690_ _0739_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_117_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4360_ _2231_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3311_ _0515_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4291_ GCDdpath0.B_reg\[95\] net251 _2170_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3242_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__buf_2
X_3173_ _1222_ _0939_ _0921_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2957_ _1003_ _1007_ _0900_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_162_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2888_ net357 GCDdpath0.B_reg\[72\] VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _2414_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_170_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4558_ _2313_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3509_ _1012_ _1527_ _0878_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4489_ GCDdpath0.B_reg\[37\] net187 _2314_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput140 operands_bits_B[10] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xinput151 operands_bits_B[11] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_1
Xinput162 operands_bits_B[14] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_1
Xinput173 operands_bits_B[24] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_2
Xinput184 operands_bits_B[34] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_1
Xinput195 operands_bits_B[44] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_127_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3860_ _1354_ _1820_ _1830_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2811_ _0855_ _0858_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__or3b_1
XFILLER_0_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3791_ _0732_ _0735_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_171_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2742_ GCDdpath0.B_reg\[39\] net320 VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2673_ _0719_ _0722_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_132_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4412_ _2267_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4343_ GCDdpath0.B_reg\[80\] net235 _2213_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4274_ _2141_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3225_ _0807_ _1259_ net390 _1212_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__and4b_1
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3156_ _0774_ _0777_ _0776_ _0772_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_145_Left_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3087_ GCDdpath0.B_reg\[120\] net283 VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3989_ _0641_ _1939_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3010_ _1056_ _1057_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4961_ clknet_leaf_34_clk _0293_ _0037_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3912_ net320 _1793_ _1873_ _0573_ _1874_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4892_ _2457_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3843_ _1806_ _1814_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3774_ _0840_ _1464_ _0571_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2725_ GCDdpath0.B_reg\[45\] net327 VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_933 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2656_ _0652_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_977 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2587_ _0607_ _0634_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4326_ GCDdpath0.B_reg\[85\] net240 _2199_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__mux2_1
X_4257_ net267 _2157_ _2158_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3208_ _1117_ _1258_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__nor2_1
X_4188_ net289 _2109_ _1282_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3139_ _0711_ _1188_ _1189_ _0841_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_174_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_162_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_166_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2510_ _0558_ _0559_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3490_ _1343_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5160_ clknet_leaf_6_clk _0492_ _0236_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_166_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4111_ _0630_ _2016_ _0620_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__a21o_1
X_5091_ clknet_leaf_32_clk _0423_ _0167_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4042_ net300 _1985_ _1911_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4944_ clknet_leaf_44_clk _0276_ _0020_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4875_ _2455_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3826_ _0737_ _1771_ _0733_ VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_691 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3757_ _0725_ _0726_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2708_ _0731_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3688_ net356 _1349_ _1681_ _1682_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2639_ _0685_ _0689_ _0672_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__a21o_1
Xoutput263 net263 VGND VGND VPWR VPWR result_bits_data[102] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput274 net274 VGND VGND VPWR VPWR result_bits_data[112] sky130_fd_sc_hd__clkbuf_4
Xoutput285 net285 VGND VGND VPWR VPWR result_bits_data[122] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput296 net296 VGND VGND VPWR VPWR result_bits_data[17] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4309_ GCDdpath0.B_reg\[90\] net246 _2184_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_163_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2990_ _1039_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_173_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4660_ _2420_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3611_ net367 net108 _1615_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4591_ _2393_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3542_ net378 _1445_ _1555_ _1556_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3473_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5143_ clknet_leaf_17_clk _0475_ _0219_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dfrtp_4
X_5074_ clknet_leaf_42_clk _0406_ _0150_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4025_ _1971_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4927_ clknet_leaf_0_clk _0259_ _0003_ VGND VGND VPWR VPWR GCDdpath0.B_reg\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4858_ _2447_ VGND VGND VPWR VPWR _2452_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_43_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3809_ GCDdpath0.B_reg\[53\] _1437_ _1300_ _1785_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__o22a_1
X_4789_ _2441_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_171_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_164_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_170_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_163_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_159_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_1045 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2973_ net266 GCDdpath0.B_reg\[105\] VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4712_ _2428_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4643_ _2413_ VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4574_ _2381_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3525_ GCDdpath0.B_reg\[93\] _1437_ _1343_ _1541_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3456_ _1318_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3387_ _1420_ _1421_ _1080_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__a21boi_2
X_5126_ clknet_leaf_15_clk _0458_ _0202_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dfrtp_4
X_5057_ clknet_leaf_39_clk _0389_ _0133_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4008_ _1938_ _1955_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_45_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_4 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3310_ _1353_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__buf_2
XFILLER_0_120_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4290_ _2181_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3241_ _1291_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__clkbuf_4
X_3172_ GCDdpath0.B_reg\[74\] net359 VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__and2b_1
XFILLER_0_174_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_174_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_961 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2956_ _1004_ _1006_ _0906_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_161_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2887_ _0934_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_161_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4626_ _2414_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_1005 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4557_ _2369_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3508_ _0998_ _1526_ _0911_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__a21o_1
X_4488_ _2321_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3439_ _1464_ _1447_ _1465_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_55_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ clknet_leaf_25_clk _0441_ _0185_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_161_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput130 operands_bits_B[100] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_1
Xinput141 operands_bits_B[110] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xinput152 operands_bits_B[120] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xinput163 operands_bits_B[15] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_1
Xinput174 operands_bits_B[25] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_2
Xinput185 operands_bits_B[35] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
Xinput196 operands_bits_B[45] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2810_ _0859_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3790_ _1769_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _0782_ _0785_ _0788_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__or4_2
XFILLER_0_125_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2672_ net347 GCDdpath0.B_reg\[63\] VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_132_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4411_ net344 _2266_ _2258_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4342_ _2218_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4273_ _2169_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__clkbuf_1
X_3224_ _1106_ _1261_ _1258_ net389 _1274_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__o41a_1
.ends

