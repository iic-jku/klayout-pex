.SUBCKT cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5
CAP1 C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5
.ENDS cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5
