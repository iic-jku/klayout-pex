* Extracted by KLayout with SKY130 LVS runset on : 11/10/2024 20:14

.SUBCKT sidewall_non_parallel_li1
.ENDS sidewall_non_parallel_li1
