* NGSPICE file created from r_wire_voltage_divider_li1.ext - technology: sky130A

.subckt r_wire_voltage_divider_li1 B A C
R0 A C.n0 426.668
R1 C.n0 B 413.868
R2 C.n0 C 72.5338
R3 A.n0 A 426.668
R4 B A.n0 413.868
R5 A.n0 C 72.5338
R6 A B.n0 426.668
R7 B.n0 B 413.868
R8 B.n0 C 72.5338
C0 B VSUBS 0.968643f
.ends
